magic
tech sky130A
magscale 1 2
timestamp 1608157713
<< locali >>
rect 22109 15351 22143 15657
rect 29377 12835 29411 12937
rect 26617 12087 26651 12257
rect 23397 11611 23431 11781
rect 41797 11067 41831 11169
rect 45017 7735 45051 7837
rect 16313 7191 16347 7293
rect 37565 5763 37599 5865
rect 43729 5559 43763 5729
rect 54585 5151 54619 5321
rect 11621 4607 11655 4777
rect 35081 4471 35115 4777
<< viali >>
rect 14381 17289 14415 17323
rect 19901 17289 19935 17323
rect 25605 17289 25639 17323
rect 40049 17289 40083 17323
rect 45569 17289 45603 17323
rect 12817 17153 12851 17187
rect 37381 17153 37415 17187
rect 13093 17085 13127 17119
rect 16957 17085 16991 17119
rect 18337 17085 18371 17119
rect 18613 17085 18647 17119
rect 22753 17085 22787 17119
rect 24041 17085 24075 17119
rect 24317 17085 24351 17119
rect 28089 17085 28123 17119
rect 34161 17085 34195 17119
rect 35633 17085 35667 17119
rect 37013 17085 37047 17119
rect 38485 17085 38519 17119
rect 38761 17085 38795 17119
rect 44005 17085 44039 17119
rect 44281 17085 44315 17119
rect 48421 17085 48455 17119
rect 49893 17085 49927 17119
rect 16773 17017 16807 17051
rect 22569 17017 22603 17051
rect 27905 17017 27939 17051
rect 33977 17017 34011 17051
rect 35449 17017 35483 17051
rect 36001 17017 36035 17051
rect 36829 17017 36863 17051
rect 48237 17017 48271 17051
rect 49709 17017 49743 17051
rect 17049 16949 17083 16983
rect 22845 16949 22879 16983
rect 28181 16949 28215 16983
rect 34253 16949 34287 16983
rect 48513 16949 48547 16983
rect 49985 16949 50019 16983
rect 18061 16745 18095 16779
rect 24133 16745 24167 16779
rect 33793 16745 33827 16779
rect 39221 16745 39255 16779
rect 47225 16745 47259 16779
rect 50813 16745 50847 16779
rect 13461 16677 13495 16711
rect 15301 16677 15335 16711
rect 19165 16677 19199 16711
rect 21373 16677 21407 16711
rect 29377 16677 29411 16711
rect 30205 16677 30239 16711
rect 40325 16677 40359 16711
rect 56977 16677 57011 16711
rect 11805 16609 11839 16643
rect 12081 16609 12115 16643
rect 15485 16609 15519 16643
rect 16681 16609 16715 16643
rect 16957 16609 16991 16643
rect 19349 16609 19383 16643
rect 21557 16609 21591 16643
rect 27721 16609 27755 16643
rect 30389 16609 30423 16643
rect 32689 16609 32723 16643
rect 35173 16609 35207 16643
rect 37841 16609 37875 16643
rect 38117 16609 38151 16643
rect 40509 16609 40543 16643
rect 43361 16609 43395 16643
rect 45845 16609 45879 16643
rect 49433 16609 49467 16643
rect 55321 16609 55355 16643
rect 55597 16609 55631 16643
rect 15853 16541 15887 16575
rect 22753 16541 22787 16575
rect 23029 16541 23063 16575
rect 27997 16541 28031 16575
rect 32413 16541 32447 16575
rect 34897 16541 34931 16575
rect 36277 16541 36311 16575
rect 43637 16541 43671 16575
rect 46121 16541 46155 16575
rect 49709 16541 49743 16575
rect 19441 16405 19475 16439
rect 21649 16405 21683 16439
rect 30481 16405 30515 16439
rect 40601 16405 40635 16439
rect 44741 16405 44775 16439
rect 13093 16201 13127 16235
rect 18521 16201 18555 16235
rect 22017 16201 22051 16235
rect 25237 16201 25271 16235
rect 30849 16201 30883 16235
rect 33885 16201 33919 16235
rect 37657 16201 37691 16235
rect 39221 16201 39255 16235
rect 44741 16201 44775 16235
rect 49433 16201 49467 16235
rect 12633 16133 12667 16167
rect 16221 16133 16255 16167
rect 18061 16133 18095 16167
rect 27261 16133 27295 16167
rect 41981 16133 42015 16167
rect 22753 16065 22787 16099
rect 23949 16065 23983 16099
rect 27997 16065 28031 16099
rect 36277 16065 36311 16099
rect 12909 15997 12943 16031
rect 14381 15997 14415 16031
rect 16497 15997 16531 16031
rect 18245 15997 18279 16031
rect 18337 15997 18371 16031
rect 20637 15997 20671 16031
rect 20729 15997 20763 16031
rect 22293 15997 22327 16031
rect 23673 15997 23707 16031
rect 27537 15997 27571 16031
rect 29285 15997 29319 16031
rect 29561 15997 29595 16031
rect 33701 15997 33735 16031
rect 34897 15997 34931 16031
rect 35081 15997 35115 16031
rect 36553 15997 36587 16031
rect 38761 15997 38795 16031
rect 38945 15997 38979 16031
rect 39037 15997 39071 16031
rect 41797 15997 41831 16031
rect 42901 15997 42935 16031
rect 43085 15997 43119 16031
rect 44281 15997 44315 16031
rect 44557 15997 44591 16031
rect 46121 15997 46155 16031
rect 46305 15997 46339 16031
rect 48053 15997 48087 16031
rect 48329 15997 48363 16031
rect 55781 15997 55815 16031
rect 12817 15929 12851 15963
rect 14197 15929 14231 15963
rect 16405 15929 16439 15963
rect 16957 15929 16991 15963
rect 21189 15929 21223 15963
rect 22201 15929 22235 15963
rect 27445 15929 27479 15963
rect 35449 15929 35483 15963
rect 43453 15929 43487 15963
rect 44465 15929 44499 15963
rect 55597 15929 55631 15963
rect 14473 15861 14507 15895
rect 46397 15861 46431 15895
rect 55873 15861 55907 15895
rect 22109 15657 22143 15691
rect 7481 15589 7515 15623
rect 12265 15589 12299 15623
rect 14197 15589 14231 15623
rect 18613 15589 18647 15623
rect 5549 15521 5583 15555
rect 5733 15521 5767 15555
rect 7665 15521 7699 15555
rect 10885 15521 10919 15555
rect 12173 15521 12207 15555
rect 12357 15521 12391 15555
rect 13645 15521 13679 15555
rect 13829 15521 13863 15555
rect 15485 15521 15519 15555
rect 16957 15521 16991 15555
rect 17233 15521 17267 15555
rect 19441 15521 19475 15555
rect 15669 15385 15703 15419
rect 22201 15589 22235 15623
rect 24961 15589 24995 15623
rect 28733 15589 28767 15623
rect 29285 15589 29319 15623
rect 36277 15589 36311 15623
rect 38485 15589 38519 15623
rect 43637 15589 43671 15623
rect 45201 15589 45235 15623
rect 45753 15589 45787 15623
rect 47501 15589 47535 15623
rect 48053 15589 48087 15623
rect 49157 15589 49191 15623
rect 49709 15589 49743 15623
rect 22845 15521 22879 15555
rect 23213 15521 23247 15555
rect 24409 15521 24443 15555
rect 24501 15521 24535 15555
rect 27077 15521 27111 15555
rect 28825 15521 28859 15555
rect 30941 15521 30975 15555
rect 36369 15521 36403 15555
rect 38393 15521 38427 15555
rect 38577 15521 38611 15555
rect 43729 15521 43763 15555
rect 45293 15521 45327 15555
rect 47593 15521 47627 15555
rect 49249 15521 49283 15555
rect 50997 15521 51031 15555
rect 51181 15521 51215 15555
rect 52377 15521 52411 15555
rect 52561 15521 52595 15555
rect 55873 15521 55907 15555
rect 56057 15521 56091 15555
rect 22753 15453 22787 15487
rect 23305 15453 23339 15487
rect 32873 15453 32907 15487
rect 33149 15453 33183 15487
rect 36093 15453 36127 15487
rect 51549 15453 51583 15487
rect 52929 15453 52963 15487
rect 24225 15385 24259 15419
rect 27261 15385 27295 15419
rect 28549 15385 28583 15419
rect 43453 15385 43487 15419
rect 5825 15317 5859 15351
rect 7757 15317 7791 15351
rect 11069 15317 11103 15351
rect 12541 15317 12575 15351
rect 19625 15317 19659 15351
rect 22109 15317 22143 15351
rect 31125 15317 31159 15351
rect 34253 15317 34287 15351
rect 36553 15317 36587 15351
rect 38761 15317 38795 15351
rect 43913 15317 43947 15351
rect 45017 15317 45051 15351
rect 47317 15317 47351 15351
rect 48973 15317 49007 15351
rect 56149 15317 56183 15351
rect 8585 15113 8619 15147
rect 15393 15113 15427 15147
rect 16313 15113 16347 15147
rect 16773 15113 16807 15147
rect 24133 15113 24167 15147
rect 25513 15113 25547 15147
rect 27997 15113 28031 15147
rect 33701 15113 33735 15147
rect 35633 15113 35667 15147
rect 39037 15113 39071 15147
rect 43545 15113 43579 15147
rect 44741 15113 44775 15147
rect 47685 15113 47719 15147
rect 53297 15113 53331 15147
rect 55413 15113 55447 15147
rect 13829 14977 13863 15011
rect 23673 14977 23707 15011
rect 35173 14977 35207 15011
rect 37381 14977 37415 15011
rect 51733 14977 51767 15011
rect 5365 14909 5399 14943
rect 5549 14909 5583 14943
rect 7021 14909 7055 14943
rect 7297 14909 7331 14943
rect 11161 14909 11195 14943
rect 12449 14909 12483 14943
rect 12725 14909 12759 14943
rect 15209 14909 15243 14943
rect 16497 14909 16531 14943
rect 16589 14909 16623 14943
rect 18521 14909 18555 14943
rect 18797 14909 18831 14943
rect 22201 14909 22235 14943
rect 22293 14909 22327 14943
rect 22569 14909 22603 14943
rect 22661 14909 22695 14943
rect 23949 14909 23983 14943
rect 25421 14909 25455 14943
rect 26801 14909 26835 14943
rect 27813 14909 27847 14943
rect 30941 14909 30975 14943
rect 32137 14909 32171 14943
rect 33333 14909 33367 14943
rect 33517 14909 33551 14943
rect 35357 14909 35391 14943
rect 35449 14909 35483 14943
rect 37473 14909 37507 14943
rect 37841 14909 37875 14943
rect 38025 14909 38059 14943
rect 38853 14909 38887 14943
rect 43361 14909 43395 14943
rect 44649 14909 44683 14943
rect 46305 14909 46339 14943
rect 47501 14909 47535 14943
rect 52009 14909 52043 14943
rect 55045 14909 55079 14943
rect 55229 14909 55263 14943
rect 10977 14841 11011 14875
rect 11529 14841 11563 14875
rect 21557 14841 21591 14875
rect 23857 14841 23891 14875
rect 25237 14841 25271 14875
rect 30757 14841 30791 14875
rect 33425 14841 33459 14875
rect 36829 14841 36863 14875
rect 44465 14841 44499 14875
rect 46121 14841 46155 14875
rect 55137 14841 55171 14875
rect 5641 14773 5675 14807
rect 19901 14773 19935 14807
rect 26893 14773 26927 14807
rect 31033 14773 31067 14807
rect 32321 14773 32355 14807
rect 46397 14773 46431 14807
rect 6009 14569 6043 14603
rect 8493 14569 8527 14603
rect 15485 14569 15519 14603
rect 43821 14569 43855 14603
rect 51641 14569 51675 14603
rect 10333 14501 10367 14535
rect 18337 14501 18371 14535
rect 21649 14501 21683 14535
rect 23673 14501 23707 14535
rect 28825 14501 28859 14535
rect 32965 14501 32999 14535
rect 33517 14501 33551 14535
rect 34529 14501 34563 14535
rect 35909 14501 35943 14535
rect 39037 14501 39071 14535
rect 46397 14501 46431 14535
rect 52929 14501 52963 14535
rect 53481 14501 53515 14535
rect 56241 14501 56275 14535
rect 58725 14501 58759 14535
rect 4629 14433 4663 14467
rect 7113 14433 7147 14467
rect 10517 14433 10551 14467
rect 15301 14433 15335 14467
rect 16681 14433 16715 14467
rect 19441 14433 19475 14467
rect 19533 14433 19567 14467
rect 19993 14433 20027 14467
rect 22293 14433 22327 14467
rect 22661 14433 22695 14467
rect 24317 14433 24351 14467
rect 24685 14433 24719 14467
rect 26709 14433 26743 14467
rect 26893 14433 26927 14467
rect 29469 14433 29503 14467
rect 29561 14433 29595 14467
rect 29837 14433 29871 14467
rect 30849 14433 30883 14467
rect 33149 14433 33183 14467
rect 34621 14433 34655 14467
rect 36093 14433 36127 14467
rect 37921 14433 37955 14467
rect 39681 14433 39715 14467
rect 40049 14433 40083 14467
rect 43637 14433 43671 14467
rect 44741 14433 44775 14467
rect 47225 14433 47259 14467
rect 50261 14433 50295 14467
rect 53021 14433 53055 14467
rect 54585 14433 54619 14467
rect 4905 14365 4939 14399
rect 7389 14365 7423 14399
rect 11713 14365 11747 14399
rect 11989 14365 12023 14399
rect 13093 14365 13127 14399
rect 16957 14365 16991 14399
rect 22385 14365 22419 14399
rect 22753 14365 22787 14399
rect 24409 14365 24443 14399
rect 24777 14365 24811 14399
rect 29929 14365 29963 14399
rect 39589 14365 39623 14399
rect 40141 14365 40175 14399
rect 45017 14365 45051 14399
rect 50537 14365 50571 14399
rect 54861 14365 54895 14399
rect 57069 14365 57103 14399
rect 57345 14365 57379 14399
rect 31033 14297 31067 14331
rect 34345 14297 34379 14331
rect 38117 14297 38151 14331
rect 10609 14229 10643 14263
rect 26985 14229 27019 14263
rect 34805 14229 34839 14263
rect 36185 14229 36219 14263
rect 47409 14229 47443 14263
rect 52745 14229 52779 14263
rect 6837 14025 6871 14059
rect 12449 14025 12483 14059
rect 12909 14025 12943 14059
rect 14473 14025 14507 14059
rect 18429 14025 18463 14059
rect 22477 14025 22511 14059
rect 24593 14025 24627 14059
rect 32965 14025 32999 14059
rect 35081 14025 35115 14059
rect 44097 14025 44131 14059
rect 46121 14025 46155 14059
rect 46581 14025 46615 14059
rect 52193 14025 52227 14059
rect 53757 14025 53791 14059
rect 55321 14025 55355 14059
rect 48053 13957 48087 13991
rect 50721 13957 50755 13991
rect 51733 13957 51767 13991
rect 5917 13889 5951 13923
rect 7573 13889 7607 13923
rect 14013 13889 14047 13923
rect 18153 13889 18187 13923
rect 19533 13889 19567 13923
rect 25881 13889 25915 13923
rect 27261 13889 27295 13923
rect 30205 13889 30239 13923
rect 31585 13889 31619 13923
rect 32689 13889 32723 13923
rect 36921 13889 36955 13923
rect 54493 13889 54527 13923
rect 56057 13889 56091 13923
rect 5273 13821 5307 13855
rect 5365 13821 5399 13855
rect 5457 13821 5491 13855
rect 7021 13821 7055 13855
rect 7113 13821 7147 13855
rect 10977 13821 11011 13855
rect 11069 13821 11103 13855
rect 11345 13821 11379 13855
rect 11529 13821 11563 13855
rect 12725 13821 12759 13855
rect 14289 13821 14323 13855
rect 18245 13821 18279 13855
rect 19809 13821 19843 13855
rect 22109 13821 22143 13855
rect 22293 13821 22327 13855
rect 24317 13821 24351 13855
rect 24409 13821 24443 13855
rect 26157 13821 26191 13855
rect 30481 13821 30515 13855
rect 32781 13821 32815 13855
rect 34897 13821 34931 13855
rect 36829 13821 36863 13855
rect 37197 13821 37231 13855
rect 37381 13821 37415 13855
rect 38853 13821 38887 13855
rect 38945 13821 38979 13855
rect 39221 13821 39255 13855
rect 39405 13821 39439 13855
rect 44649 13821 44683 13855
rect 44741 13821 44775 13855
rect 45017 13821 45051 13855
rect 45201 13821 45235 13855
rect 46397 13821 46431 13855
rect 47869 13821 47903 13855
rect 48973 13821 49007 13855
rect 50537 13821 50571 13855
rect 51917 13821 51951 13855
rect 52009 13821 52043 13855
rect 54033 13821 54067 13855
rect 55505 13821 55539 13855
rect 55597 13821 55631 13855
rect 10333 13753 10367 13787
rect 12633 13753 12667 13787
rect 14197 13753 14231 13787
rect 22201 13753 22235 13787
rect 36185 13753 36219 13787
rect 38209 13753 38243 13787
rect 46305 13753 46339 13787
rect 53941 13753 53975 13787
rect 21097 13685 21131 13719
rect 49157 13685 49191 13719
rect 25513 13481 25547 13515
rect 42901 13481 42935 13515
rect 54953 13481 54987 13515
rect 5365 13413 5399 13447
rect 10425 13413 10459 13447
rect 11437 13413 11471 13447
rect 17141 13413 17175 13447
rect 18981 13413 19015 13447
rect 20913 13413 20947 13447
rect 26525 13413 26559 13447
rect 28365 13413 28399 13447
rect 32321 13413 32355 13447
rect 33885 13413 33919 13447
rect 36645 13413 36679 13447
rect 37749 13413 37783 13447
rect 41521 13413 41555 13447
rect 44557 13413 44591 13447
rect 48973 13413 49007 13447
rect 52469 13413 52503 13447
rect 54677 13413 54711 13447
rect 5273 13345 5307 13379
rect 5457 13345 5491 13379
rect 9781 13345 9815 13379
rect 10149 13345 10183 13379
rect 12081 13345 12115 13379
rect 12449 13345 12483 13379
rect 13553 13345 13587 13379
rect 15301 13345 15335 13379
rect 17601 13345 17635 13379
rect 17969 13345 18003 13379
rect 19441 13345 19475 13379
rect 19809 13345 19843 13379
rect 21373 13345 21407 13379
rect 21557 13345 21591 13379
rect 21741 13345 21775 13379
rect 22753 13345 22787 13379
rect 22845 13345 22879 13379
rect 24133 13345 24167 13379
rect 25329 13345 25363 13379
rect 27077 13345 27111 13379
rect 27353 13345 27387 13379
rect 28549 13345 28583 13379
rect 30389 13345 30423 13379
rect 30573 13345 30607 13379
rect 30757 13345 30791 13379
rect 32413 13345 32447 13379
rect 33977 13345 34011 13379
rect 36185 13345 36219 13379
rect 38393 13345 38427 13379
rect 38485 13345 38519 13379
rect 38761 13345 38795 13379
rect 38945 13345 38979 13379
rect 41705 13345 41739 13379
rect 43085 13345 43119 13379
rect 45201 13345 45235 13379
rect 45569 13345 45603 13379
rect 46765 13345 46799 13379
rect 47501 13345 47535 13379
rect 47869 13345 47903 13379
rect 48053 13345 48087 13379
rect 49617 13345 49651 13379
rect 49985 13345 50019 13379
rect 51181 13345 51215 13379
rect 53113 13345 53147 13379
rect 53447 13345 53481 13379
rect 54861 13345 54895 13379
rect 11989 13277 12023 13311
rect 12541 13277 12575 13311
rect 13461 13277 13495 13311
rect 18061 13277 18095 13311
rect 19901 13277 19935 13311
rect 27537 13277 27571 13311
rect 36093 13277 36127 13311
rect 45109 13277 45143 13311
rect 45661 13277 45695 13311
rect 47409 13277 47443 13311
rect 49525 13277 49559 13311
rect 50077 13277 50111 13311
rect 51089 13277 51123 13311
rect 51641 13277 51675 13311
rect 53205 13277 53239 13311
rect 53573 13277 53607 13311
rect 15485 13209 15519 13243
rect 30205 13209 30239 13243
rect 46949 13209 46983 13243
rect 5641 13141 5675 13175
rect 13737 13141 13771 13175
rect 23029 13141 23063 13175
rect 24317 13141 24351 13175
rect 28641 13141 28675 13175
rect 32137 13141 32171 13175
rect 32597 13141 32631 13175
rect 33701 13141 33735 13175
rect 34161 13141 34195 13175
rect 41797 13141 41831 13175
rect 46581 13141 46615 13175
rect 4813 12937 4847 12971
rect 10425 12937 10459 12971
rect 18245 12937 18279 12971
rect 22293 12937 22327 12971
rect 29377 12937 29411 12971
rect 29653 12937 29687 12971
rect 32045 12937 32079 12971
rect 40785 12937 40819 12971
rect 45201 12937 45235 12971
rect 46213 12937 46247 12971
rect 50537 12937 50571 12971
rect 52745 12937 52779 12971
rect 54769 12937 54803 12971
rect 23857 12869 23891 12903
rect 25881 12869 25915 12903
rect 48329 12869 48363 12903
rect 6837 12801 6871 12835
rect 7389 12801 7423 12835
rect 13001 12801 13035 12835
rect 13553 12801 13587 12835
rect 19809 12801 19843 12835
rect 20545 12801 20579 12835
rect 21833 12801 21867 12835
rect 29377 12801 29411 12835
rect 32689 12801 32723 12835
rect 36645 12801 36679 12835
rect 40509 12801 40543 12835
rect 42533 12801 42567 12835
rect 43361 12801 43395 12835
rect 43913 12801 43947 12835
rect 46857 12801 46891 12835
rect 47225 12801 47259 12835
rect 53205 12801 53239 12835
rect 53757 12801 53791 12835
rect 55229 12801 55263 12835
rect 58357 12801 58391 12835
rect 5365 12733 5399 12767
rect 5457 12733 5491 12767
rect 5733 12733 5767 12767
rect 5917 12733 5951 12767
rect 6929 12733 6963 12767
rect 9229 12733 9263 12767
rect 10977 12733 11011 12767
rect 11069 12733 11103 12767
rect 11345 12733 11379 12767
rect 11529 12733 11563 12767
rect 13093 12733 13127 12767
rect 13461 12733 13495 12767
rect 14473 12733 14507 12767
rect 15761 12733 15795 12767
rect 16589 12733 16623 12767
rect 16773 12733 16807 12767
rect 18429 12733 18463 12767
rect 18521 12733 18555 12767
rect 20453 12733 20487 12767
rect 20821 12733 20855 12767
rect 20913 12733 20947 12767
rect 22109 12733 22143 12767
rect 23673 12733 23707 12767
rect 26065 12733 26099 12767
rect 26433 12733 26467 12767
rect 26525 12733 26559 12767
rect 27629 12733 27663 12767
rect 29469 12733 29503 12767
rect 30757 12733 30791 12767
rect 32597 12733 32631 12767
rect 32965 12733 32999 12767
rect 33057 12733 33091 12767
rect 34989 12733 35023 12767
rect 36093 12733 36127 12767
rect 36205 12733 36239 12767
rect 37473 12733 37507 12767
rect 37585 12733 37619 12767
rect 38025 12733 38059 12767
rect 40601 12733 40635 12767
rect 41981 12733 42015 12767
rect 42073 12733 42107 12767
rect 44189 12733 44223 12767
rect 44373 12733 44407 12767
rect 45385 12733 45419 12767
rect 46765 12733 46799 12767
rect 47133 12733 47167 12767
rect 48145 12733 48179 12767
rect 50261 12733 50295 12767
rect 50353 12733 50387 12767
rect 53297 12733 53331 12767
rect 53665 12733 53699 12767
rect 55321 12733 55355 12767
rect 55689 12733 55723 12767
rect 55781 12733 55815 12767
rect 58633 12733 58667 12767
rect 12449 12665 12483 12699
rect 17141 12665 17175 12699
rect 18981 12665 19015 12699
rect 22017 12665 22051 12699
rect 27445 12665 27479 12699
rect 30573 12665 30607 12699
rect 9413 12597 9447 12631
rect 14657 12597 14691 12631
rect 15577 12597 15611 12631
rect 27721 12597 27755 12631
rect 30849 12597 30883 12631
rect 35173 12597 35207 12631
rect 59737 12597 59771 12631
rect 9965 12393 9999 12427
rect 23029 12393 23063 12427
rect 24317 12393 24351 12427
rect 30665 12393 30699 12427
rect 49985 12393 50019 12427
rect 5365 12325 5399 12359
rect 7941 12325 7975 12359
rect 17417 12325 17451 12359
rect 18981 12325 19015 12359
rect 30757 12325 30791 12359
rect 31125 12325 31159 12359
rect 32137 12325 32171 12359
rect 36645 12325 36679 12359
rect 44557 12325 44591 12359
rect 47133 12325 47167 12359
rect 52469 12325 52503 12359
rect 54585 12325 54619 12359
rect 6009 12257 6043 12291
rect 6377 12257 6411 12291
rect 6561 12257 6595 12291
rect 7481 12257 7515 12291
rect 9781 12257 9815 12291
rect 11529 12257 11563 12291
rect 11897 12257 11931 12291
rect 11989 12257 12023 12291
rect 13001 12257 13035 12291
rect 16037 12257 16071 12291
rect 16221 12257 16255 12291
rect 17601 12257 17635 12291
rect 19809 12257 19843 12291
rect 19993 12257 20027 12291
rect 21741 12257 21775 12291
rect 22753 12257 22787 12291
rect 22937 12257 22971 12291
rect 24133 12257 24167 12291
rect 25329 12257 25363 12291
rect 26617 12257 26651 12291
rect 26709 12257 26743 12291
rect 26893 12257 26927 12291
rect 27261 12257 27295 12291
rect 28549 12257 28583 12291
rect 28733 12257 28767 12291
rect 28917 12257 28951 12291
rect 29377 12257 29411 12291
rect 29561 12257 29595 12291
rect 30573 12257 30607 12291
rect 32781 12257 32815 12291
rect 33115 12257 33149 12291
rect 33333 12257 33367 12291
rect 34345 12257 34379 12291
rect 34437 12257 34471 12291
rect 36185 12257 36219 12291
rect 41245 12257 41279 12291
rect 41705 12257 41739 12291
rect 42073 12257 42107 12291
rect 43361 12257 43395 12291
rect 45201 12257 45235 12291
rect 45569 12257 45603 12291
rect 45753 12257 45787 12291
rect 46673 12257 46707 12291
rect 49801 12257 49835 12291
rect 50905 12257 50939 12291
rect 50997 12257 51031 12291
rect 53113 12257 53147 12291
rect 53481 12257 53515 12291
rect 53665 12257 53699 12291
rect 55229 12257 55263 12291
rect 55597 12257 55631 12291
rect 55781 12257 55815 12291
rect 58173 12257 58207 12291
rect 58357 12257 58391 12291
rect 58541 12257 58575 12291
rect 5917 12189 5951 12223
rect 7389 12189 7423 12223
rect 10885 12189 10919 12223
rect 11437 12189 11471 12223
rect 12909 12189 12943 12223
rect 16589 12189 16623 12223
rect 17969 12189 18003 12223
rect 19533 12189 19567 12223
rect 20913 12189 20947 12223
rect 21465 12189 21499 12223
rect 21925 12189 21959 12223
rect 28089 12189 28123 12223
rect 30389 12189 30423 12223
rect 32873 12189 32907 12223
rect 36093 12189 36127 12223
rect 38761 12189 38795 12223
rect 39037 12189 39071 12223
rect 42165 12189 42199 12223
rect 45109 12189 45143 12223
rect 46581 12189 46615 12223
rect 51457 12189 51491 12223
rect 53021 12189 53055 12223
rect 55137 12189 55171 12223
rect 34161 12121 34195 12155
rect 43545 12121 43579 12155
rect 57989 12121 58023 12155
rect 13185 12053 13219 12087
rect 25513 12053 25547 12087
rect 26617 12053 26651 12087
rect 34621 12053 34655 12087
rect 40141 12053 40175 12087
rect 6929 11849 6963 11883
rect 20085 11849 20119 11883
rect 22293 11849 22327 11883
rect 35173 11849 35207 11883
rect 46397 11849 46431 11883
rect 12541 11781 12575 11815
rect 23397 11781 23431 11815
rect 23857 11781 23891 11815
rect 48605 11781 48639 11815
rect 52009 11781 52043 11815
rect 3065 11713 3099 11747
rect 7573 11713 7607 11747
rect 7941 11713 7975 11747
rect 11529 11713 11563 11747
rect 13001 11713 13035 11747
rect 13553 11713 13587 11747
rect 15393 11713 15427 11747
rect 18429 11713 18463 11747
rect 21097 11713 21131 11747
rect 3157 11645 3191 11679
rect 4445 11645 4479 11679
rect 4905 11645 4939 11679
rect 5089 11645 5123 11679
rect 5365 11645 5399 11679
rect 5549 11645 5583 11679
rect 5917 11645 5951 11679
rect 7481 11645 7515 11679
rect 7849 11645 7883 11679
rect 8861 11645 8895 11679
rect 9045 11645 9079 11679
rect 10977 11645 11011 11679
rect 11069 11645 11103 11679
rect 13093 11645 13127 11679
rect 13461 11645 13495 11679
rect 14933 11645 14967 11679
rect 15301 11645 15335 11679
rect 16497 11645 16531 11679
rect 16773 11645 16807 11679
rect 17141 11645 17175 11679
rect 18705 11645 18739 11679
rect 20637 11645 20671 11679
rect 20729 11645 20763 11679
rect 21005 11645 21039 11679
rect 22201 11645 22235 11679
rect 26893 11713 26927 11747
rect 28089 11713 28123 11747
rect 30573 11713 30607 11747
rect 31585 11713 31619 11747
rect 32137 11713 32171 11747
rect 32597 11713 32631 11747
rect 33977 11713 34011 11747
rect 41889 11713 41923 11747
rect 44097 11713 44131 11747
rect 45109 11713 45143 11747
rect 46121 11713 46155 11747
rect 52653 11713 52687 11747
rect 54309 11713 54343 11747
rect 57989 11713 58023 11747
rect 23673 11645 23707 11679
rect 24777 11645 24811 11679
rect 25881 11645 25915 11679
rect 27445 11645 27479 11679
rect 27537 11645 27571 11679
rect 27721 11645 27755 11679
rect 28273 11645 28307 11679
rect 30205 11645 30239 11679
rect 32413 11645 32447 11679
rect 33609 11645 33643 11679
rect 35081 11645 35115 11679
rect 36369 11645 36403 11679
rect 36645 11645 36679 11679
rect 41613 11645 41647 11679
rect 44649 11645 44683 11679
rect 44925 11645 44959 11679
rect 46213 11645 46247 11679
rect 48789 11645 48823 11679
rect 49157 11645 49191 11679
rect 49249 11645 49283 11679
rect 50537 11645 50571 11679
rect 52193 11645 52227 11679
rect 52561 11645 52595 11679
rect 53757 11645 53791 11679
rect 53849 11645 53883 11679
rect 55873 11645 55907 11679
rect 56241 11645 56275 11679
rect 56333 11645 56367 11679
rect 57713 11645 57747 11679
rect 3617 11577 3651 11611
rect 14473 11577 14507 11611
rect 16589 11577 16623 11611
rect 18797 11577 18831 11611
rect 19165 11577 19199 11611
rect 22017 11577 22051 11611
rect 23397 11577 23431 11611
rect 30021 11577 30055 11611
rect 33425 11577 33459 11611
rect 34897 11577 34931 11611
rect 55413 11577 55447 11611
rect 9137 11509 9171 11543
rect 16313 11509 16347 11543
rect 18613 11509 18647 11543
rect 24961 11509 24995 11543
rect 25973 11509 26007 11543
rect 37749 11509 37783 11543
rect 43177 11509 43211 11543
rect 50721 11509 50755 11543
rect 59093 11509 59127 11543
rect 24409 11305 24443 11339
rect 28457 11305 28491 11339
rect 29837 11305 29871 11339
rect 31125 11305 31159 11339
rect 32321 11305 32355 11339
rect 40601 11305 40635 11339
rect 53113 11305 53147 11339
rect 57989 11305 58023 11339
rect 59093 11305 59127 11339
rect 3157 11237 3191 11271
rect 6929 11237 6963 11271
rect 11345 11237 11379 11271
rect 15853 11237 15887 11271
rect 17325 11237 17359 11271
rect 18705 11237 18739 11271
rect 21465 11237 21499 11271
rect 26801 11237 26835 11271
rect 28181 11237 28215 11271
rect 29561 11237 29595 11271
rect 44189 11237 44223 11271
rect 48053 11237 48087 11271
rect 50629 11237 50663 11271
rect 55137 11237 55171 11271
rect 2605 11169 2639 11203
rect 2789 11169 2823 11203
rect 4445 11169 4479 11203
rect 7481 11169 7515 11203
rect 7757 11169 7791 11203
rect 7941 11169 7975 11203
rect 9689 11169 9723 11203
rect 10793 11169 10827 11203
rect 10885 11169 10919 11203
rect 15301 11169 15335 11203
rect 15393 11169 15427 11203
rect 17509 11169 17543 11203
rect 19349 11169 19383 11203
rect 19717 11169 19751 11203
rect 19809 11169 19843 11203
rect 21005 11169 21039 11203
rect 22569 11169 22603 11203
rect 23121 11169 23155 11203
rect 23305 11169 23339 11203
rect 24225 11169 24259 11203
rect 25329 11169 25363 11203
rect 26893 11169 26927 11203
rect 28365 11169 28399 11203
rect 29745 11169 29779 11203
rect 30941 11169 30975 11203
rect 32137 11169 32171 11203
rect 34897 11169 34931 11203
rect 36277 11169 36311 11203
rect 36645 11169 36679 11203
rect 37755 11169 37789 11203
rect 41797 11169 41831 11203
rect 41889 11169 41923 11203
rect 42073 11169 42107 11203
rect 42441 11169 42475 11203
rect 43637 11169 43671 11203
rect 43729 11169 43763 11203
rect 47593 11169 47627 11203
rect 48973 11169 49007 11203
rect 49249 11169 49283 11203
rect 52009 11169 52043 11203
rect 54677 11169 54711 11203
rect 56425 11169 56459 11203
rect 56701 11169 56735 11203
rect 58909 11169 58943 11203
rect 4721 11101 4755 11135
rect 12173 11101 12207 11135
rect 12449 11101 12483 11135
rect 17877 11101 17911 11135
rect 19441 11101 19475 11135
rect 20913 11101 20947 11135
rect 33241 11101 33275 11135
rect 33517 11101 33551 11135
rect 36737 11101 36771 11135
rect 39221 11101 39255 11135
rect 39497 11101 39531 11135
rect 45017 11101 45051 11135
rect 45293 11101 45327 11135
rect 47501 11101 47535 11135
rect 51733 11101 51767 11135
rect 54585 11101 54619 11135
rect 5825 11033 5859 11067
rect 9873 11033 9907 11067
rect 13737 11033 13771 11067
rect 25513 11033 25547 11067
rect 36093 11033 36127 11067
rect 37933 11033 37967 11067
rect 41797 11033 41831 11067
rect 23397 10965 23431 10999
rect 26617 10965 26651 10999
rect 27077 10965 27111 10999
rect 46397 10965 46431 10999
rect 7113 10761 7147 10795
rect 8953 10761 8987 10795
rect 18797 10761 18831 10795
rect 36277 10761 36311 10795
rect 43729 10761 43763 10795
rect 49893 10761 49927 10795
rect 53205 10761 53239 10795
rect 14105 10693 14139 10727
rect 16405 10693 16439 10727
rect 19073 10693 19107 10727
rect 33241 10693 33275 10727
rect 38485 10693 38519 10727
rect 55689 10693 55723 10727
rect 3249 10625 3283 10659
rect 12541 10625 12575 10659
rect 12817 10625 12851 10659
rect 19809 10625 19843 10659
rect 21097 10625 21131 10659
rect 22753 10625 22787 10659
rect 25237 10625 25271 10659
rect 26617 10625 26651 10659
rect 26893 10625 26927 10659
rect 29745 10625 29779 10659
rect 35173 10625 35207 10659
rect 42165 10625 42199 10659
rect 45109 10625 45143 10659
rect 46121 10625 46155 10659
rect 48329 10625 48363 10659
rect 57345 10625 57379 10659
rect 2881 10557 2915 10591
rect 4077 10557 4111 10591
rect 4353 10557 4387 10591
rect 6837 10557 6871 10591
rect 6929 10557 6963 10591
rect 8769 10557 8803 10591
rect 9873 10557 9907 10591
rect 10977 10557 11011 10591
rect 11069 10557 11103 10591
rect 15025 10557 15059 10591
rect 15301 10557 15335 10591
rect 18981 10557 19015 10591
rect 19349 10557 19383 10591
rect 20821 10557 20855 10591
rect 21373 10557 21407 10591
rect 23673 10557 23707 10591
rect 25329 10557 25363 10591
rect 28273 10557 28307 10591
rect 29469 10557 29503 10591
rect 30665 10557 30699 10591
rect 31861 10557 31895 10591
rect 33425 10557 33459 10591
rect 33609 10557 33643 10591
rect 33769 10557 33803 10591
rect 34897 10557 34931 10591
rect 38669 10557 38703 10591
rect 38853 10557 38887 10591
rect 39037 10557 39071 10591
rect 42441 10557 42475 10591
rect 44833 10557 44867 10591
rect 46581 10557 46615 10591
rect 46949 10557 46983 10591
rect 47041 10557 47075 10591
rect 48605 10557 48639 10591
rect 51733 10557 51767 10591
rect 52929 10557 52963 10591
rect 53021 10557 53055 10591
rect 54309 10557 54343 10591
rect 55873 10557 55907 10591
rect 56057 10557 56091 10591
rect 56241 10557 56275 10591
rect 57621 10557 57655 10591
rect 2697 10489 2731 10523
rect 11529 10489 11563 10523
rect 19257 10489 19291 10523
rect 25789 10489 25823 10523
rect 29285 10489 29319 10523
rect 44649 10489 44683 10523
rect 5641 10421 5675 10455
rect 10057 10421 10091 10455
rect 20637 10421 20671 10455
rect 23857 10421 23891 10455
rect 30849 10421 30883 10455
rect 32045 10421 32079 10455
rect 51825 10421 51859 10455
rect 54493 10421 54527 10455
rect 58725 10421 58759 10455
rect 5641 10217 5675 10251
rect 34989 10217 35023 10251
rect 36369 10217 36403 10251
rect 47041 10217 47075 10251
rect 7113 10149 7147 10183
rect 11437 10149 11471 10183
rect 15301 10149 15335 10183
rect 19533 10149 19567 10183
rect 19625 10149 19659 10183
rect 23857 10149 23891 10183
rect 25605 10149 25639 10183
rect 28825 10149 28859 10183
rect 36093 10149 36127 10183
rect 39405 10149 39439 10183
rect 48973 10149 49007 10183
rect 55781 10149 55815 10183
rect 6653 10081 6687 10115
rect 10057 10081 10091 10115
rect 12081 10081 12115 10115
rect 12449 10081 12483 10115
rect 12633 10081 12667 10115
rect 13461 10081 13495 10115
rect 15761 10081 15795 10115
rect 15945 10081 15979 10115
rect 16129 10081 16163 10115
rect 17969 10081 18003 10115
rect 19441 10081 19475 10115
rect 21097 10081 21131 10115
rect 22201 10081 22235 10115
rect 22477 10081 22511 10115
rect 25053 10081 25087 10115
rect 25145 10081 25179 10115
rect 26801 10081 26835 10115
rect 27077 10081 27111 10115
rect 27537 10081 27571 10115
rect 27721 10081 27755 10115
rect 29009 10081 29043 10115
rect 30205 10081 30239 10115
rect 32321 10081 32355 10115
rect 33609 10081 33643 10115
rect 36277 10081 36311 10115
rect 37749 10081 37783 10115
rect 39865 10081 39899 10115
rect 40049 10081 40083 10115
rect 40233 10081 40267 10115
rect 41705 10081 41739 10115
rect 42073 10081 42107 10115
rect 42165 10081 42199 10115
rect 44373 10081 44407 10115
rect 46029 10081 46063 10115
rect 46857 10081 46891 10115
rect 49433 10081 49467 10115
rect 49801 10081 49835 10115
rect 54677 10081 54711 10115
rect 56241 10081 56275 10115
rect 56609 10081 56643 10115
rect 4077 10013 4111 10047
rect 4353 10013 4387 10047
rect 6561 10013 6595 10047
rect 9965 10013 9999 10047
rect 11989 10013 12023 10047
rect 13829 10013 13863 10047
rect 17877 10013 17911 10047
rect 19257 10013 19291 10047
rect 19993 10013 20027 10047
rect 32229 10013 32263 10047
rect 32781 10013 32815 10047
rect 33885 10013 33919 10047
rect 44649 10013 44683 10047
rect 49893 10013 49927 10047
rect 51549 10013 51583 10047
rect 51825 10013 51859 10047
rect 56701 10013 56735 10047
rect 57621 10013 57655 10047
rect 57897 10013 57931 10047
rect 21281 9945 21315 9979
rect 26617 9945 26651 9979
rect 30389 9945 30423 9979
rect 41521 9945 41555 9979
rect 10241 9877 10275 9911
rect 13599 9877 13633 9911
rect 13737 9877 13771 9911
rect 14105 9877 14139 9911
rect 18153 9877 18187 9911
rect 29101 9877 29135 9911
rect 37933 9877 37967 9911
rect 53113 9877 53147 9911
rect 54861 9877 54895 9911
rect 59001 9877 59035 9911
rect 10241 9673 10275 9707
rect 37013 9673 37047 9707
rect 44419 9673 44453 9707
rect 44557 9673 44591 9707
rect 49065 9673 49099 9707
rect 7113 9605 7147 9639
rect 15209 9605 15243 9639
rect 17049 9605 17083 9639
rect 23765 9605 23799 9639
rect 33241 9605 33275 9639
rect 50077 9605 50111 9639
rect 2973 9537 3007 9571
rect 12449 9537 12483 9571
rect 15853 9537 15887 9571
rect 18889 9537 18923 9571
rect 22753 9537 22787 9571
rect 26709 9537 26743 9571
rect 29745 9537 29779 9571
rect 39589 9537 39623 9571
rect 43453 9537 43487 9571
rect 44649 9537 44683 9571
rect 46121 9537 46155 9571
rect 48237 9537 48271 9571
rect 59461 9537 59495 9571
rect 3249 9469 3283 9503
rect 7297 9469 7331 9503
rect 7481 9469 7515 9503
rect 7665 9469 7699 9503
rect 8677 9469 8711 9503
rect 8953 9469 8987 9503
rect 11161 9469 11195 9503
rect 12725 9469 12759 9503
rect 15393 9469 15427 9503
rect 15761 9469 15795 9503
rect 16865 9469 16899 9503
rect 18337 9469 18371 9503
rect 18429 9469 18463 9503
rect 19717 9469 19751 9503
rect 19993 9469 20027 9503
rect 22201 9469 22235 9503
rect 22293 9469 22327 9503
rect 23673 9469 23707 9503
rect 25329 9469 25363 9503
rect 25513 9469 25547 9503
rect 25881 9469 25915 9503
rect 27261 9469 27295 9503
rect 27445 9469 27479 9503
rect 27629 9469 27663 9503
rect 27813 9469 27847 9503
rect 28181 9469 28215 9503
rect 29469 9469 29503 9503
rect 32597 9469 32631 9503
rect 33425 9469 33459 9503
rect 33793 9469 33827 9503
rect 33885 9469 33919 9503
rect 35357 9469 35391 9503
rect 35541 9469 35575 9503
rect 35725 9469 35759 9503
rect 36737 9469 36771 9503
rect 36829 9469 36863 9503
rect 39037 9469 39071 9503
rect 39129 9469 39163 9503
rect 41429 9469 41463 9503
rect 41797 9469 41831 9503
rect 42073 9469 42107 9503
rect 46397 9469 46431 9503
rect 47685 9469 47719 9503
rect 47777 9469 47811 9503
rect 49249 9469 49283 9503
rect 50261 9469 50295 9503
rect 50445 9469 50479 9503
rect 50629 9469 50663 9503
rect 52653 9469 52687 9503
rect 52929 9469 52963 9503
rect 55413 9469 55447 9503
rect 58081 9469 58115 9503
rect 58357 9469 58391 9503
rect 14105 9401 14139 9435
rect 21373 9401 21407 9435
rect 29285 9401 29319 9435
rect 30757 9401 30791 9435
rect 34897 9401 34931 9435
rect 44281 9401 44315 9435
rect 46489 9401 46523 9435
rect 46857 9401 46891 9435
rect 55229 9401 55263 9435
rect 55781 9401 55815 9435
rect 4353 9333 4387 9367
rect 11345 9333 11379 9367
rect 32045 9333 32079 9367
rect 32781 9333 32815 9367
rect 41245 9333 41279 9367
rect 44925 9333 44959 9367
rect 46305 9333 46339 9367
rect 54033 9333 54067 9367
rect 2145 9061 2179 9095
rect 4721 9061 4755 9095
rect 17049 9061 17083 9095
rect 20913 9061 20947 9095
rect 23305 9061 23339 9095
rect 24869 9061 24903 9095
rect 28733 9061 28767 9095
rect 35633 9061 35667 9095
rect 38301 9061 38335 9095
rect 41797 9061 41831 9095
rect 46397 9061 46431 9095
rect 46581 9061 46615 9095
rect 49433 9061 49467 9095
rect 50813 9061 50847 9095
rect 56057 9061 56091 9095
rect 58081 9061 58115 9095
rect 2605 8993 2639 9027
rect 2973 8993 3007 9027
rect 5181 8993 5215 9027
rect 5549 8993 5583 9027
rect 5641 8993 5675 9027
rect 8309 8993 8343 9027
rect 10333 8993 10367 9027
rect 10701 8993 10735 9027
rect 12357 8993 12391 9027
rect 12725 8993 12759 9027
rect 12909 8993 12943 9027
rect 13737 8993 13771 9027
rect 13921 8993 13955 9027
rect 16221 8993 16255 9027
rect 16589 8993 16623 9027
rect 17969 8993 18003 9027
rect 19257 8993 19291 9027
rect 19404 8993 19438 9027
rect 21557 8993 21591 9027
rect 21925 8993 21959 9027
rect 23121 8993 23155 9027
rect 23213 8993 23247 9027
rect 24777 8993 24811 9027
rect 30021 8993 30055 9027
rect 30665 8993 30699 9027
rect 32137 8993 32171 9027
rect 34805 8993 34839 9027
rect 36093 8993 36127 9027
rect 36461 8993 36495 9027
rect 36553 8993 36587 9027
rect 37841 8993 37875 9027
rect 39865 8993 39899 9027
rect 40049 8993 40083 9027
rect 41337 8993 41371 9027
rect 44189 8993 44223 9027
rect 44741 8993 44775 9027
rect 44925 8993 44959 9027
rect 46489 8993 46523 9027
rect 47961 8993 47995 9027
rect 49617 8993 49651 9027
rect 49985 8993 50019 9027
rect 51457 8993 51491 9027
rect 51825 8993 51859 9027
rect 51917 8993 51951 9027
rect 52837 8993 52871 9027
rect 54769 8993 54803 9027
rect 56701 8993 56735 9027
rect 57069 8993 57103 9027
rect 57253 8993 57287 9027
rect 58725 8993 58759 9027
rect 59093 8993 59127 9027
rect 60197 8993 60231 9027
rect 60289 8993 60323 9027
rect 3065 8925 3099 8959
rect 8217 8925 8251 8959
rect 8769 8925 8803 8959
rect 10241 8925 10275 8959
rect 10793 8925 10827 8959
rect 11713 8925 11747 8959
rect 12265 8925 12299 8959
rect 16497 8925 16531 8959
rect 17877 8925 17911 8959
rect 18429 8925 18463 8959
rect 19625 8925 19659 8959
rect 21465 8925 21499 8959
rect 22017 8925 22051 8959
rect 22937 8925 22971 8959
rect 23673 8925 23707 8959
rect 27077 8925 27111 8959
rect 27353 8925 27387 8959
rect 32229 8925 32263 8959
rect 33149 8925 33183 8959
rect 33425 8925 33459 8959
rect 37749 8925 37783 8959
rect 41245 8925 41279 8959
rect 44005 8925 44039 8959
rect 46213 8925 46247 8959
rect 46949 8925 46983 8959
rect 51365 8925 51399 8959
rect 52984 8925 53018 8959
rect 53205 8925 53239 8959
rect 54677 8925 54711 8959
rect 56793 8925 56827 8959
rect 58817 8925 58851 8959
rect 59185 8925 59219 8959
rect 45109 8857 45143 8891
rect 53297 8857 53331 8891
rect 9781 8789 9815 8823
rect 14013 8789 14047 8823
rect 16037 8789 16071 8823
rect 19533 8789 19567 8823
rect 19901 8789 19935 8823
rect 30205 8789 30239 8823
rect 30849 8789 30883 8823
rect 40141 8789 40175 8823
rect 47777 8789 47811 8823
rect 53113 8789 53147 8823
rect 54953 8789 54987 8823
rect 60473 8789 60507 8823
rect 1961 8585 1995 8619
rect 4261 8585 4295 8619
rect 5549 8585 5583 8619
rect 9689 8585 9723 8619
rect 21097 8585 21131 8619
rect 37105 8585 37139 8619
rect 38393 8585 38427 8619
rect 39497 8585 39531 8619
rect 41705 8585 41739 8619
rect 43729 8585 43763 8619
rect 50537 8585 50571 8619
rect 52745 8585 52779 8619
rect 13553 8517 13587 8551
rect 23857 8517 23891 8551
rect 46213 8517 46247 8551
rect 58817 8517 58851 8551
rect 2881 8449 2915 8483
rect 8401 8449 8435 8483
rect 12909 8449 12943 8483
rect 14749 8449 14783 8483
rect 15945 8449 15979 8483
rect 22569 8449 22603 8483
rect 25697 8449 25731 8483
rect 26709 8449 26743 8483
rect 30205 8449 30239 8483
rect 31861 8449 31895 8483
rect 32413 8449 32447 8483
rect 33609 8449 33643 8483
rect 46949 8449 46983 8483
rect 53297 8449 53331 8483
rect 55045 8449 55079 8483
rect 55137 8449 55171 8483
rect 1869 8381 1903 8415
rect 3157 8381 3191 8415
rect 5365 8381 5399 8415
rect 8125 8381 8159 8415
rect 10609 8381 10643 8415
rect 10977 8381 11011 8415
rect 11161 8381 11195 8415
rect 13277 8381 13311 8415
rect 13645 8381 13679 8415
rect 14657 8381 14691 8415
rect 16037 8381 16071 8415
rect 18521 8381 18555 8415
rect 18705 8381 18739 8415
rect 19073 8381 19107 8415
rect 19901 8381 19935 8415
rect 20085 8381 20119 8415
rect 20545 8381 20579 8415
rect 20637 8381 20671 8415
rect 22293 8381 22327 8415
rect 23673 8381 23707 8415
rect 25237 8381 25271 8415
rect 25421 8381 25455 8415
rect 26985 8381 27019 8415
rect 27353 8381 27387 8415
rect 29653 8381 29687 8415
rect 29745 8381 29779 8415
rect 31953 8381 31987 8415
rect 33241 8381 33275 8415
rect 33793 8381 33827 8415
rect 34897 8381 34931 8415
rect 35449 8381 35483 8415
rect 35725 8381 35759 8415
rect 36829 8381 36863 8415
rect 36921 8381 36955 8415
rect 38209 8381 38243 8415
rect 39313 8381 39347 8415
rect 40509 8381 40543 8415
rect 42257 8381 42291 8415
rect 42349 8381 42383 8415
rect 42625 8381 42659 8415
rect 42809 8381 42843 8415
rect 44203 8381 44237 8415
rect 44373 8381 44407 8415
rect 44649 8381 44683 8415
rect 44833 8381 44867 8415
rect 45845 8381 45879 8415
rect 46305 8381 46339 8415
rect 46857 8381 46891 8415
rect 48237 8381 48271 8415
rect 50261 8381 50295 8415
rect 50353 8381 50387 8415
rect 53219 8381 53253 8415
rect 53665 8381 53699 8415
rect 53849 8381 53883 8415
rect 55873 8381 55907 8415
rect 56011 8381 56045 8415
rect 58541 8381 58575 8415
rect 59277 8381 59311 8415
rect 59553 8381 59587 8415
rect 16497 8313 16531 8347
rect 22109 8313 22143 8347
rect 27629 8313 27663 8347
rect 36001 8313 36035 8347
rect 48053 8313 48087 8347
rect 40693 8245 40727 8279
rect 45661 8245 45695 8279
rect 48329 8245 48363 8279
rect 9965 8041 9999 8075
rect 46489 8041 46523 8075
rect 47777 8041 47811 8075
rect 55229 8041 55263 8075
rect 56609 8041 56643 8075
rect 4261 7973 4295 8007
rect 8217 7973 8251 8007
rect 12081 7973 12115 8007
rect 26801 7973 26835 8007
rect 33885 7973 33919 8007
rect 39589 7973 39623 8007
rect 58541 7973 58575 8007
rect 2605 7905 2639 7939
rect 2973 7905 3007 7939
rect 4721 7905 4755 7939
rect 5089 7905 5123 7939
rect 5181 7905 5215 7939
rect 8401 7905 8435 7939
rect 10333 7905 10367 7939
rect 10701 7905 10735 7939
rect 10885 7905 10919 7939
rect 11989 7905 12023 7939
rect 12541 7905 12575 7939
rect 12909 7905 12943 7939
rect 14105 7905 14139 7939
rect 15393 7905 15427 7939
rect 17601 7905 17635 7939
rect 17785 7905 17819 7939
rect 19533 7905 19567 7939
rect 19809 7905 19843 7939
rect 20913 7905 20947 7939
rect 21097 7905 21131 7939
rect 22477 7905 22511 7939
rect 23029 7905 23063 7939
rect 27467 7905 27501 7939
rect 27813 7905 27847 7939
rect 27997 7905 28031 7939
rect 29009 7905 29043 7939
rect 29101 7905 29135 7939
rect 30665 7905 30699 7939
rect 31125 7905 31159 7939
rect 32597 7905 32631 7939
rect 34529 7905 34563 7939
rect 34897 7905 34931 7939
rect 34989 7905 35023 7939
rect 36001 7905 36035 7939
rect 36093 7905 36127 7939
rect 36226 7905 36260 7939
rect 37749 7905 37783 7939
rect 39129 7905 39163 7939
rect 40417 7905 40451 7939
rect 41153 7905 41187 7939
rect 41981 7905 42015 7939
rect 43637 7905 43671 7939
rect 44097 7905 44131 7939
rect 47593 7905 47627 7939
rect 51089 7905 51123 7939
rect 51457 7905 51491 7939
rect 53205 7905 53239 7939
rect 54769 7905 54803 7939
rect 55045 7905 55079 7939
rect 56793 7905 56827 7939
rect 56977 7905 57011 7939
rect 57345 7905 57379 7939
rect 58633 7905 58667 7939
rect 60289 7905 60323 7939
rect 3065 7837 3099 7871
rect 8769 7837 8803 7871
rect 10241 7837 10275 7871
rect 13001 7837 13035 7871
rect 15301 7837 15335 7871
rect 16773 7837 16807 7871
rect 17325 7837 17359 7871
rect 18981 7837 19015 7871
rect 19993 7837 20027 7871
rect 21373 7837 21407 7871
rect 23121 7837 23155 7871
rect 27353 7837 27387 7871
rect 32505 7837 32539 7871
rect 34437 7837 34471 7871
rect 36645 7837 36679 7871
rect 39037 7837 39071 7871
rect 45017 7837 45051 7871
rect 45109 7837 45143 7871
rect 45385 7837 45419 7871
rect 50813 7837 50847 7871
rect 53113 7837 53147 7871
rect 53665 7837 53699 7871
rect 57253 7837 57287 7871
rect 60197 7837 60231 7871
rect 2421 7769 2455 7803
rect 22569 7769 22603 7803
rect 30481 7769 30515 7803
rect 42165 7769 42199 7803
rect 51457 7769 51491 7803
rect 54861 7769 54895 7803
rect 11805 7701 11839 7735
rect 14289 7701 14323 7735
rect 15577 7701 15611 7735
rect 28825 7701 28859 7735
rect 29285 7701 29319 7735
rect 32781 7701 32815 7735
rect 37933 7701 37967 7735
rect 40509 7701 40543 7735
rect 43453 7701 43487 7735
rect 45017 7701 45051 7735
rect 58357 7701 58391 7735
rect 58817 7701 58851 7735
rect 60473 7701 60507 7735
rect 5641 7497 5675 7531
rect 12725 7497 12759 7531
rect 16405 7497 16439 7531
rect 19901 7497 19935 7531
rect 25789 7429 25823 7463
rect 27169 7429 27203 7463
rect 31953 7429 31987 7463
rect 2881 7361 2915 7395
rect 5365 7361 5399 7395
rect 8309 7361 8343 7395
rect 15025 7361 15059 7395
rect 17141 7361 17175 7395
rect 21005 7361 21039 7395
rect 21557 7361 21591 7395
rect 33609 7361 33643 7395
rect 41337 7361 41371 7395
rect 44189 7361 44223 7395
rect 44741 7361 44775 7395
rect 47133 7361 47167 7395
rect 56057 7361 56091 7395
rect 58541 7361 58575 7395
rect 3157 7293 3191 7327
rect 5457 7293 5491 7327
rect 8585 7293 8619 7327
rect 10793 7293 10827 7327
rect 10885 7293 10919 7327
rect 11069 7293 11103 7327
rect 12909 7293 12943 7327
rect 13093 7293 13127 7327
rect 13461 7293 13495 7327
rect 13645 7293 13679 7327
rect 14473 7293 14507 7327
rect 14606 7293 14640 7327
rect 16221 7293 16255 7327
rect 16313 7293 16347 7327
rect 16722 7293 16756 7327
rect 18521 7293 18555 7327
rect 18797 7293 18831 7327
rect 21833 7293 21867 7327
rect 22017 7293 22051 7327
rect 24225 7293 24259 7327
rect 24317 7293 24351 7327
rect 25605 7293 25639 7327
rect 27353 7293 27387 7327
rect 27721 7293 27755 7327
rect 27813 7293 27847 7327
rect 29469 7293 29503 7327
rect 30665 7293 30699 7327
rect 31769 7293 31803 7327
rect 33241 7293 33275 7327
rect 33977 7293 34011 7327
rect 35541 7293 35575 7327
rect 36093 7293 36127 7327
rect 36277 7293 36311 7327
rect 36645 7293 36679 7327
rect 37013 7293 37047 7327
rect 39221 7293 39255 7327
rect 39589 7293 39623 7327
rect 41245 7293 41279 7327
rect 42073 7293 42107 7327
rect 42165 7293 42199 7327
rect 43085 7293 43119 7327
rect 45017 7293 45051 7327
rect 45201 7293 45235 7327
rect 46673 7293 46707 7327
rect 46949 7293 46983 7327
rect 48697 7293 48731 7327
rect 50537 7293 50571 7327
rect 52285 7293 52319 7327
rect 52561 7293 52595 7327
rect 55781 7293 55815 7327
rect 56241 7293 56275 7327
rect 57345 7293 57379 7327
rect 58817 7293 58851 7327
rect 9965 7225 9999 7259
rect 11529 7225 11563 7259
rect 16589 7225 16623 7259
rect 24777 7225 24811 7259
rect 29285 7225 29319 7259
rect 35725 7225 35759 7259
rect 39034 7225 39068 7259
rect 46121 7225 46155 7259
rect 53941 7225 53975 7259
rect 4445 7157 4479 7191
rect 16037 7157 16071 7191
rect 16313 7157 16347 7191
rect 29561 7157 29595 7191
rect 30849 7157 30883 7191
rect 43269 7157 43303 7191
rect 48881 7157 48915 7191
rect 50721 7157 50755 7191
rect 57529 7157 57563 7191
rect 59921 7157 59955 7191
rect 3065 6953 3099 6987
rect 34253 6953 34287 6987
rect 37841 6953 37875 6987
rect 45661 6953 45695 6987
rect 17693 6885 17727 6919
rect 18705 6885 18739 6919
rect 27169 6885 27203 6919
rect 52469 6885 52503 6919
rect 58081 6885 58115 6919
rect 60749 6885 60783 6919
rect 2973 6817 3007 6851
rect 4077 6817 4111 6851
rect 5733 6817 5767 6851
rect 6653 6817 6687 6851
rect 8217 6817 8251 6851
rect 8585 6817 8619 6851
rect 9689 6817 9723 6851
rect 10609 6817 10643 6851
rect 11897 6817 11931 6851
rect 12587 6817 12621 6851
rect 12725 6817 12759 6851
rect 13829 6817 13863 6851
rect 14013 6817 14047 6851
rect 19349 6817 19383 6851
rect 19717 6817 19751 6851
rect 20913 6817 20947 6851
rect 21465 6817 21499 6851
rect 22937 6817 22971 6851
rect 23397 6817 23431 6851
rect 25053 6817 25087 6851
rect 25237 6817 25271 6851
rect 25421 6817 25455 6851
rect 26985 6817 27019 6851
rect 27537 6817 27571 6851
rect 27997 6817 28031 6851
rect 28089 6817 28123 6851
rect 28457 6817 28491 6851
rect 29837 6817 29871 6851
rect 30941 6817 30975 6851
rect 32689 6817 32723 6851
rect 33793 6817 33827 6851
rect 34069 6817 34103 6851
rect 35817 6817 35851 6851
rect 36001 6817 36035 6851
rect 36185 6817 36219 6851
rect 36369 6817 36403 6851
rect 36645 6817 36679 6851
rect 37749 6817 37783 6851
rect 38761 6817 38795 6851
rect 38945 6817 38979 6851
rect 39313 6817 39347 6851
rect 40325 6817 40359 6851
rect 40417 6817 40451 6851
rect 40877 6817 40911 6851
rect 41889 6817 41923 6851
rect 41981 6817 42015 6851
rect 43361 6817 43395 6851
rect 43913 6817 43947 6851
rect 44189 6817 44223 6851
rect 45201 6817 45235 6851
rect 45477 6817 45511 6851
rect 46765 6817 46799 6851
rect 47041 6817 47075 6851
rect 49065 6817 49099 6851
rect 51089 6817 51123 6851
rect 51181 6817 51215 6851
rect 53113 6817 53147 6851
rect 53481 6817 53515 6851
rect 54769 6817 54803 6851
rect 54953 6817 54987 6851
rect 56701 6817 56735 6851
rect 56977 6817 57011 6851
rect 57253 6817 57287 6851
rect 58725 6817 58759 6851
rect 58817 6817 58851 6851
rect 59093 6817 59127 6851
rect 60289 6817 60323 6851
rect 4353 6749 4387 6783
rect 6561 6749 6595 6783
rect 8401 6749 8435 6783
rect 10701 6749 10735 6783
rect 11989 6749 12023 6783
rect 16037 6749 16071 6783
rect 16313 6749 16347 6783
rect 19257 6749 19291 6783
rect 19809 6749 19843 6783
rect 22845 6749 22879 6783
rect 35357 6749 35391 6783
rect 40141 6749 40175 6783
rect 41705 6749 41739 6783
rect 42441 6749 42475 6783
rect 44373 6749 44407 6783
rect 47317 6749 47351 6783
rect 48973 6749 49007 6783
rect 49525 6749 49559 6783
rect 53205 6749 53239 6783
rect 53573 6749 53607 6783
rect 55321 6749 55355 6783
rect 56241 6749 56275 6783
rect 59185 6749 59219 6783
rect 60197 6749 60231 6783
rect 10149 6681 10183 6715
rect 21005 6681 21039 6715
rect 24869 6681 24903 6715
rect 31125 6681 31159 6715
rect 32873 6681 32907 6715
rect 33885 6681 33919 6715
rect 45293 6681 45327 6715
rect 46857 6681 46891 6715
rect 6837 6613 6871 6647
rect 14105 6613 14139 6647
rect 30021 6613 30055 6647
rect 51365 6613 51399 6647
rect 9689 6409 9723 6443
rect 28181 6409 28215 6443
rect 40785 6409 40819 6443
rect 53297 6409 53331 6443
rect 16497 6341 16531 6375
rect 21373 6341 21407 6375
rect 52101 6341 52135 6375
rect 53665 6341 53699 6375
rect 3709 6273 3743 6307
rect 10149 6273 10183 6307
rect 10701 6273 10735 6307
rect 12449 6273 12483 6307
rect 16957 6273 16991 6307
rect 19533 6273 19567 6307
rect 25237 6273 25271 6307
rect 31447 6273 31481 6307
rect 39037 6273 39071 6307
rect 39589 6273 39623 6307
rect 47961 6273 47995 6307
rect 50261 6273 50295 6307
rect 53389 6273 53423 6307
rect 60105 6273 60139 6307
rect 2697 6205 2731 6239
rect 4169 6205 4203 6239
rect 4537 6205 4571 6239
rect 4629 6205 4663 6239
rect 7021 6205 7055 6239
rect 8217 6205 8251 6239
rect 10241 6205 10275 6239
rect 10609 6205 10643 6239
rect 13185 6205 13219 6239
rect 15209 6205 15243 6239
rect 16405 6205 16439 6239
rect 16681 6205 16715 6239
rect 18061 6205 18095 6239
rect 19441 6205 19475 6239
rect 20269 6205 20303 6239
rect 20361 6205 20395 6239
rect 21281 6205 21315 6239
rect 21557 6205 21591 6239
rect 23857 6205 23891 6239
rect 24961 6205 24995 6239
rect 27997 6205 28031 6239
rect 29285 6205 29319 6239
rect 31309 6205 31343 6239
rect 31585 6205 31619 6239
rect 33589 6205 33623 6239
rect 34897 6205 34931 6239
rect 36185 6205 36219 6239
rect 36461 6205 36495 6239
rect 36921 6205 36955 6239
rect 37289 6205 37323 6239
rect 37749 6205 37783 6239
rect 39129 6205 39163 6239
rect 40693 6205 40727 6239
rect 41889 6205 41923 6239
rect 42625 6205 42659 6239
rect 42901 6205 42935 6239
rect 44649 6205 44683 6239
rect 44741 6205 44775 6239
rect 45201 6205 45235 6239
rect 46581 6205 46615 6239
rect 46949 6205 46983 6239
rect 47869 6205 47903 6239
rect 48697 6205 48731 6239
rect 48789 6205 48823 6239
rect 50394 6205 50428 6239
rect 51917 6205 51951 6239
rect 53168 6205 53202 6239
rect 54585 6205 54619 6239
rect 55137 6205 55171 6239
rect 55413 6205 55447 6239
rect 55597 6205 55631 6239
rect 58725 6205 58759 6239
rect 58817 6205 58851 6239
rect 59093 6205 59127 6239
rect 59185 6205 59219 6239
rect 60565 6205 60599 6239
rect 60749 6205 60783 6239
rect 60933 6205 60967 6239
rect 6837 6137 6871 6171
rect 12817 6137 12851 6171
rect 15025 6137 15059 6171
rect 30757 6137 30791 6171
rect 33425 6137 33459 6171
rect 33977 6137 34011 6171
rect 36369 6137 36403 6171
rect 40509 6137 40543 6171
rect 46397 6137 46431 6171
rect 50813 6137 50847 6171
rect 53021 6137 53055 6171
rect 58081 6137 58115 6171
rect 2789 6069 2823 6103
rect 7113 6069 7147 6103
rect 8309 6069 8343 6103
rect 12633 6069 12667 6103
rect 12725 6069 12759 6103
rect 15301 6069 15335 6103
rect 18245 6069 18279 6103
rect 21741 6069 21775 6103
rect 24041 6069 24075 6103
rect 26525 6069 26559 6103
rect 29469 6069 29503 6103
rect 35081 6069 35115 6103
rect 41981 6069 42015 6103
rect 37565 5865 37599 5899
rect 38301 5865 38335 5899
rect 49433 5865 49467 5899
rect 53113 5865 53147 5899
rect 4169 5797 4203 5831
rect 23305 5797 23339 5831
rect 26525 5797 26559 5831
rect 32137 5797 32171 5831
rect 34897 5797 34931 5831
rect 41337 5797 41371 5831
rect 47041 5797 47075 5831
rect 49617 5797 49651 5831
rect 49985 5797 50019 5831
rect 51549 5797 51583 5831
rect 52929 5797 52963 5831
rect 53297 5797 53331 5831
rect 55321 5797 55355 5831
rect 58449 5797 58483 5831
rect 2605 5729 2639 5763
rect 2697 5729 2731 5763
rect 4629 5729 4663 5763
rect 4813 5729 4847 5763
rect 4997 5729 5031 5763
rect 6193 5729 6227 5763
rect 6561 5729 6595 5763
rect 6837 5729 6871 5763
rect 7941 5729 7975 5763
rect 8217 5729 8251 5763
rect 11069 5729 11103 5763
rect 13553 5729 13587 5763
rect 15485 5729 15519 5763
rect 15669 5729 15703 5763
rect 16865 5729 16899 5763
rect 19349 5729 19383 5763
rect 19533 5729 19567 5763
rect 23397 5729 23431 5763
rect 24869 5729 24903 5763
rect 25237 5729 25271 5763
rect 26985 5729 27019 5763
rect 27169 5729 27203 5763
rect 27445 5729 27479 5763
rect 27629 5729 27663 5763
rect 27813 5729 27847 5763
rect 28917 5729 28951 5763
rect 30987 5729 31021 5763
rect 31217 5729 31251 5763
rect 32321 5729 32355 5763
rect 34437 5729 34471 5763
rect 36461 5729 36495 5763
rect 37565 5729 37599 5763
rect 38117 5729 38151 5763
rect 39221 5729 39255 5763
rect 39405 5729 39439 5763
rect 39773 5729 39807 5763
rect 40785 5729 40819 5763
rect 40877 5729 40911 5763
rect 42165 5729 42199 5763
rect 43729 5729 43763 5763
rect 43821 5729 43855 5763
rect 44189 5729 44223 5763
rect 44465 5729 44499 5763
rect 45390 5729 45424 5763
rect 45661 5729 45695 5763
rect 47869 5729 47903 5763
rect 49525 5729 49559 5763
rect 51733 5729 51767 5763
rect 53205 5729 53239 5763
rect 56149 5729 56183 5763
rect 57161 5729 57195 5763
rect 57345 5729 57379 5763
rect 57805 5729 57839 5763
rect 57897 5729 57931 5763
rect 60197 5729 60231 5763
rect 60289 5729 60323 5763
rect 8401 5661 8435 5695
rect 11345 5661 11379 5695
rect 16037 5661 16071 5695
rect 17141 5661 17175 5695
rect 25053 5661 25087 5695
rect 28825 5661 28859 5695
rect 30205 5661 30239 5695
rect 30757 5661 30791 5695
rect 32689 5661 32723 5695
rect 34345 5661 34379 5695
rect 6929 5593 6963 5627
rect 8033 5593 8067 5627
rect 45477 5661 45511 5695
rect 46121 5661 46155 5695
rect 47593 5661 47627 5695
rect 48053 5661 48087 5695
rect 49249 5661 49283 5695
rect 53665 5661 53699 5695
rect 55873 5661 55907 5695
rect 56333 5661 56367 5695
rect 2881 5525 2915 5559
rect 12449 5525 12483 5559
rect 13737 5525 13771 5559
rect 18245 5525 18279 5559
rect 19625 5525 19659 5559
rect 23121 5525 23155 5559
rect 23581 5525 23615 5559
rect 29101 5525 29135 5559
rect 36645 5525 36679 5559
rect 40601 5525 40635 5559
rect 42349 5525 42383 5559
rect 43729 5525 43763 5559
rect 51825 5525 51859 5559
rect 60473 5525 60507 5559
rect 3065 5321 3099 5355
rect 5733 5321 5767 5355
rect 7113 5321 7147 5355
rect 12541 5321 12575 5355
rect 18061 5321 18095 5355
rect 40785 5321 40819 5355
rect 53021 5321 53055 5355
rect 54585 5321 54619 5355
rect 57621 5321 57655 5355
rect 10609 5253 10643 5287
rect 24133 5253 24167 5287
rect 26893 5253 26927 5287
rect 30481 5253 30515 5287
rect 43453 5253 43487 5287
rect 47685 5253 47719 5287
rect 50077 5253 50111 5287
rect 52837 5253 52871 5287
rect 2789 5185 2823 5219
rect 7573 5185 7607 5219
rect 11345 5185 11379 5219
rect 13185 5185 13219 5219
rect 15301 5185 15335 5219
rect 16129 5185 16163 5219
rect 18797 5185 18831 5219
rect 19717 5185 19751 5219
rect 20085 5185 20119 5219
rect 35909 5185 35943 5219
rect 44189 5185 44223 5219
rect 46397 5185 46431 5219
rect 52929 5185 52963 5219
rect 58817 5185 58851 5219
rect 2901 5117 2935 5151
rect 4169 5117 4203 5151
rect 4445 5117 4479 5151
rect 7481 5117 7515 5151
rect 7849 5117 7883 5151
rect 8033 5117 8067 5151
rect 9045 5117 9079 5151
rect 10885 5117 10919 5151
rect 13093 5117 13127 5151
rect 13461 5117 13495 5151
rect 13553 5117 13587 5151
rect 14749 5117 14783 5151
rect 14841 5117 14875 5151
rect 16681 5117 16715 5151
rect 16957 5117 16991 5151
rect 17141 5117 17175 5151
rect 18337 5117 18371 5151
rect 19625 5117 19659 5151
rect 19901 5117 19935 5151
rect 21373 5117 21407 5151
rect 24041 5117 24075 5151
rect 24501 5117 24535 5151
rect 25237 5117 25271 5151
rect 25513 5117 25547 5151
rect 25973 5117 26007 5151
rect 26801 5117 26835 5151
rect 27353 5117 27387 5151
rect 30297 5117 30331 5151
rect 31585 5117 31619 5151
rect 31953 5117 31987 5151
rect 32229 5117 32263 5151
rect 33333 5117 33367 5151
rect 34897 5117 34931 5151
rect 36461 5117 36495 5151
rect 36553 5117 36587 5151
rect 36737 5117 36771 5151
rect 36921 5117 36955 5151
rect 37289 5117 37323 5151
rect 39037 5117 39071 5151
rect 39221 5117 39255 5151
rect 39589 5117 39623 5151
rect 40693 5117 40727 5151
rect 41429 5117 41463 5151
rect 42257 5117 42291 5151
rect 43729 5117 43763 5151
rect 46121 5117 46155 5151
rect 49433 5117 49467 5151
rect 49801 5117 49835 5151
rect 50077 5117 50111 5151
rect 52708 5117 52742 5151
rect 54585 5117 54619 5151
rect 54677 5117 54711 5151
rect 54769 5117 54803 5151
rect 54953 5117 54987 5151
rect 57437 5117 57471 5151
rect 58541 5117 58575 5151
rect 8861 5049 8895 5083
rect 10793 5049 10827 5083
rect 18245 5049 18279 5083
rect 21189 5049 21223 5083
rect 43637 5049 43671 5083
rect 52561 5049 52595 5083
rect 55413 5049 55447 5083
rect 9137 4981 9171 5015
rect 21465 4981 21499 5015
rect 31493 4981 31527 5015
rect 33517 4981 33551 5015
rect 34989 4981 35023 5015
rect 42441 4981 42475 5015
rect 59921 4981 59955 5015
rect 11621 4777 11655 4811
rect 12357 4777 12391 4811
rect 28917 4777 28951 4811
rect 35081 4777 35115 4811
rect 43637 4777 43671 4811
rect 45569 4777 45603 4811
rect 3157 4709 3191 4743
rect 5365 4709 5399 4743
rect 2697 4641 2731 4675
rect 4077 4641 4111 4675
rect 5825 4641 5859 4675
rect 6193 4641 6227 4675
rect 7297 4641 7331 4675
rect 8125 4641 8159 4675
rect 8217 4641 8251 4675
rect 11713 4709 11747 4743
rect 13553 4709 13587 4743
rect 13645 4709 13679 4743
rect 15301 4709 15335 4743
rect 24133 4709 24167 4743
rect 28273 4709 28307 4743
rect 30205 4709 30239 4743
rect 13461 4641 13495 4675
rect 17693 4641 17727 4675
rect 18705 4641 18739 4675
rect 19441 4641 19475 4675
rect 22109 4641 22143 4675
rect 22477 4641 22511 4675
rect 22753 4641 22787 4675
rect 24593 4641 24627 4675
rect 24869 4641 24903 4675
rect 25053 4641 25087 4675
rect 25237 4641 25271 4675
rect 25513 4641 25547 4675
rect 26525 4641 26559 4675
rect 26617 4641 26651 4675
rect 31033 4641 31067 4675
rect 31217 4641 31251 4675
rect 32137 4641 32171 4675
rect 32413 4641 32447 4675
rect 2605 4573 2639 4607
rect 6285 4573 6319 4607
rect 7389 4573 7423 4607
rect 11621 4573 11655 4607
rect 12081 4573 12115 4607
rect 13277 4573 13311 4607
rect 14013 4573 14047 4607
rect 15669 4573 15703 4607
rect 16865 4573 16899 4607
rect 17417 4573 17451 4607
rect 17877 4573 17911 4607
rect 27077 4573 27111 4607
rect 28641 4573 28675 4607
rect 30757 4573 30791 4607
rect 18797 4505 18831 4539
rect 22201 4505 22235 4539
rect 28549 4505 28583 4539
rect 47961 4709 47995 4743
rect 50629 4709 50663 4743
rect 55781 4709 55815 4743
rect 35173 4641 35207 4675
rect 36277 4641 36311 4675
rect 36461 4641 36495 4675
rect 38393 4641 38427 4675
rect 38485 4641 38519 4675
rect 41153 4641 41187 4675
rect 41383 4641 41417 4675
rect 43361 4641 43395 4675
rect 43545 4641 43579 4675
rect 45385 4641 45419 4675
rect 46581 4641 46615 4675
rect 47869 4641 47903 4675
rect 48973 4641 49007 4675
rect 52101 4641 52135 4675
rect 52469 4641 52503 4675
rect 56379 4641 56413 4675
rect 56517 4641 56551 4675
rect 58817 4641 58851 4675
rect 36829 4573 36863 4607
rect 40601 4573 40635 4607
rect 41613 4573 41647 4607
rect 46489 4573 46523 4607
rect 47041 4573 47075 4607
rect 49249 4573 49283 4607
rect 51457 4573 51491 4607
rect 52193 4573 52227 4607
rect 52377 4573 52411 4607
rect 55689 4573 55723 4607
rect 57989 4573 58023 4607
rect 59001 4573 59035 4607
rect 35357 4505 35391 4539
rect 58449 4505 58483 4539
rect 4169 4437 4203 4471
rect 11851 4437 11885 4471
rect 11989 4437 12023 4471
rect 15439 4437 15473 4471
rect 15577 4437 15611 4471
rect 15945 4437 15979 4471
rect 28411 4437 28445 4471
rect 33701 4437 33735 4471
rect 35081 4437 35115 4471
rect 38209 4437 38243 4471
rect 38669 4437 38703 4471
rect 29929 4233 29963 4267
rect 35081 4233 35115 4267
rect 44005 4233 44039 4267
rect 49433 4165 49467 4199
rect 3157 4097 3191 4131
rect 4537 4097 4571 4131
rect 7757 4097 7791 4131
rect 18245 4097 18279 4131
rect 20177 4097 20211 4131
rect 25697 4097 25731 4131
rect 37013 4097 37047 4131
rect 39129 4097 39163 4131
rect 40601 4097 40635 4131
rect 40877 4097 40911 4131
rect 47041 4097 47075 4131
rect 52285 4097 52319 4131
rect 55505 4097 55539 4131
rect 2605 4029 2639 4063
rect 2697 4029 2731 4063
rect 3985 4029 4019 4063
rect 4077 4029 4111 4063
rect 5365 4029 5399 4063
rect 5457 4029 5491 4063
rect 5917 4029 5951 4063
rect 7297 4029 7331 4063
rect 7481 4029 7515 4063
rect 7849 4029 7883 4063
rect 8861 4029 8895 4063
rect 13093 4029 13127 4063
rect 13185 4029 13219 4063
rect 14933 4029 14967 4063
rect 15301 4029 15335 4063
rect 16681 4029 16715 4063
rect 16957 4029 16991 4063
rect 17141 4029 17175 4063
rect 18935 4029 18969 4063
rect 19061 4029 19095 4063
rect 20085 4029 20119 4063
rect 20361 4029 20395 4063
rect 22477 4029 22511 4063
rect 23765 4029 23799 4063
rect 23857 4029 23891 4063
rect 25973 4029 26007 4063
rect 26157 4029 26191 4063
rect 27169 4029 27203 4063
rect 30205 4029 30239 4063
rect 31493 4029 31527 4063
rect 31769 4029 31803 4063
rect 34897 4029 34931 4063
rect 36001 4029 36035 4063
rect 37289 4029 37323 4063
rect 39405 4029 39439 4063
rect 39589 4029 39623 4063
rect 43821 4029 43855 4063
rect 44925 4029 44959 4063
rect 47133 4029 47167 4063
rect 47501 4029 47535 4063
rect 47685 4029 47719 4063
rect 49617 4029 49651 4063
rect 49801 4029 49835 4063
rect 49985 4029 50019 4063
rect 52561 4029 52595 4063
rect 55413 4029 55447 4063
rect 55873 4029 55907 4063
rect 57437 4029 57471 4063
rect 58541 4029 58575 4063
rect 58817 4029 58851 4063
rect 13645 3961 13679 3995
rect 14749 3961 14783 3995
rect 16129 3961 16163 3995
rect 18337 3961 18371 3995
rect 24317 3961 24351 3995
rect 25145 3961 25179 3995
rect 26985 3961 27019 3995
rect 30113 3961 30147 3995
rect 30665 3961 30699 3995
rect 37197 3961 37231 3995
rect 37749 3961 37783 3995
rect 38577 3961 38611 3995
rect 46489 3961 46523 3995
rect 6929 3893 6963 3927
rect 9045 3893 9079 3927
rect 20545 3893 20579 3927
rect 22661 3893 22695 3927
rect 27261 3893 27295 3927
rect 32873 3893 32907 3927
rect 36093 3893 36127 3927
rect 41981 3893 42015 3927
rect 45109 3893 45143 3927
rect 53849 3893 53883 3927
rect 57621 3893 57655 3927
rect 59921 3893 59955 3927
rect 21097 3689 21131 3723
rect 23489 3689 23523 3723
rect 27813 3689 27847 3723
rect 32229 3689 32263 3723
rect 34345 3689 34379 3723
rect 40325 3689 40359 3723
rect 41613 3689 41647 3723
rect 49893 3689 49927 3723
rect 27721 3621 27755 3655
rect 27905 3621 27939 3655
rect 28273 3621 28307 3655
rect 29837 3621 29871 3655
rect 34529 3621 34563 3655
rect 34897 3621 34931 3655
rect 36001 3621 36035 3655
rect 36093 3621 36127 3655
rect 52929 3621 52963 3655
rect 58081 3621 58115 3655
rect 4537 3553 4571 3587
rect 6469 3553 6503 3587
rect 6837 3553 6871 3587
rect 7021 3553 7055 3587
rect 7941 3553 7975 3587
rect 8585 3553 8619 3587
rect 11989 3553 12023 3587
rect 13093 3553 13127 3587
rect 13277 3553 13311 3587
rect 16313 3553 16347 3587
rect 16497 3553 16531 3587
rect 17049 3553 17083 3587
rect 17233 3553 17267 3587
rect 18889 3553 18923 3587
rect 19349 3553 19383 3587
rect 20913 3553 20947 3587
rect 23213 3553 23247 3587
rect 23397 3553 23431 3587
rect 25421 3553 25455 3587
rect 29929 3553 29963 3587
rect 32781 3553 32815 3587
rect 33149 3553 33183 3587
rect 34437 3553 34471 3587
rect 35909 3553 35943 3587
rect 37749 3553 37783 3587
rect 39221 3553 39255 3587
rect 41429 3553 41463 3587
rect 45201 3553 45235 3587
rect 46581 3553 46615 3587
rect 49617 3553 49651 3587
rect 49801 3553 49835 3587
rect 51641 3553 51675 3587
rect 55321 3553 55355 3587
rect 55689 3553 55723 3587
rect 56793 3553 56827 3587
rect 58725 3553 58759 3587
rect 59093 3553 59127 3587
rect 59185 3553 59219 3587
rect 60197 3553 60231 3587
rect 4445 3485 4479 3519
rect 4997 3485 5031 3519
rect 6561 3485 6595 3519
rect 13645 3485 13679 3519
rect 18613 3485 18647 3519
rect 19625 3485 19659 3519
rect 24593 3485 24627 3519
rect 25145 3485 25179 3519
rect 25605 3485 25639 3519
rect 27537 3485 27571 3519
rect 29653 3485 29687 3519
rect 32597 3485 32631 3519
rect 33057 3485 33091 3519
rect 34161 3485 34195 3519
rect 35541 3485 35575 3519
rect 35725 3485 35759 3519
rect 36461 3485 36495 3519
rect 38945 3485 38979 3519
rect 46305 3485 46339 3519
rect 51549 3485 51583 3519
rect 52101 3485 52135 3519
rect 53076 3485 53110 3519
rect 53297 3485 53331 3519
rect 54677 3485 54711 3519
rect 55413 3485 55447 3519
rect 55597 3485 55631 3519
rect 56701 3485 56735 3519
rect 58633 3485 58667 3519
rect 7941 3417 7975 3451
rect 45385 3417 45419 3451
rect 5917 3349 5951 3383
rect 12173 3349 12207 3383
rect 17509 3349 17543 3383
rect 30113 3349 30147 3383
rect 37933 3349 37967 3383
rect 47869 3349 47903 3383
rect 53205 3349 53239 3383
rect 53573 3349 53607 3383
rect 56977 3349 57011 3383
rect 60289 3349 60323 3383
rect 22661 3145 22695 3179
rect 27629 3145 27663 3179
rect 39313 3145 39347 3179
rect 40674 3145 40708 3179
rect 44925 3145 44959 3179
rect 48586 3145 48620 3179
rect 52469 3145 52503 3179
rect 53481 3145 53515 3179
rect 58495 3145 58529 3179
rect 7113 3077 7147 3111
rect 14933 3077 14967 3111
rect 16037 3077 16071 3111
rect 40785 3077 40819 3111
rect 48697 3077 48731 3111
rect 58633 3077 58667 3111
rect 5273 3009 5307 3043
rect 5825 3009 5859 3043
rect 7849 3009 7883 3043
rect 13461 3009 13495 3043
rect 16589 3009 16623 3043
rect 19165 3009 19199 3043
rect 24869 3009 24903 3043
rect 28365 3009 28399 3043
rect 30481 3009 30515 3043
rect 30941 3009 30975 3043
rect 31769 3009 31803 3043
rect 32229 3009 32263 3043
rect 36461 3009 36495 3043
rect 38209 3009 38243 3043
rect 40877 3009 40911 3043
rect 41245 3009 41279 3043
rect 48789 3009 48823 3043
rect 53941 3009 53975 3043
rect 55873 3009 55907 3043
rect 58725 3009 58759 3043
rect 5365 2941 5399 2975
rect 5733 2941 5767 2975
rect 6837 2941 6871 2975
rect 7757 2941 7791 2975
rect 13369 2941 13403 2975
rect 13737 2941 13771 2975
rect 13921 2941 13955 2975
rect 14749 2941 14783 2975
rect 16511 2941 16545 2975
rect 16957 2941 16991 2975
rect 17141 2941 17175 2975
rect 18705 2941 18739 2975
rect 18797 2941 18831 2975
rect 19073 2941 19107 2975
rect 20545 2941 20579 2975
rect 20729 2941 20763 2975
rect 20913 2941 20947 2975
rect 22477 2941 22511 2975
rect 24593 2941 24627 2975
rect 27813 2941 27847 2975
rect 27905 2941 27939 2975
rect 30757 2941 30791 2975
rect 32413 2941 32447 2975
rect 32781 2941 32815 2975
rect 32965 2941 32999 2975
rect 33793 2941 33827 2975
rect 35725 2941 35759 2975
rect 37933 2941 37967 2975
rect 42073 2941 42107 2975
rect 44833 2941 44867 2975
rect 46121 2941 46155 2975
rect 46765 2941 46799 2975
rect 47041 2941 47075 2975
rect 47501 2941 47535 2975
rect 49985 2941 50019 2975
rect 52285 2941 52319 2975
rect 54033 2941 54067 2975
rect 54401 2941 54435 2975
rect 54585 2941 54619 2975
rect 55597 2941 55631 2975
rect 60105 2941 60139 2975
rect 4721 2873 4755 2907
rect 12725 2873 12759 2907
rect 18061 2873 18095 2907
rect 20085 2873 20119 2907
rect 26249 2873 26283 2907
rect 29929 2873 29963 2907
rect 36093 2873 36127 2907
rect 40509 2873 40543 2907
rect 42165 2873 42199 2907
rect 44649 2873 44683 2907
rect 48421 2873 48455 2907
rect 55413 2873 55447 2907
rect 58357 2873 58391 2907
rect 59921 2873 59955 2907
rect 33885 2805 33919 2839
rect 35909 2805 35943 2839
rect 36001 2805 36035 2839
rect 46213 2805 46247 2839
rect 49065 2805 49099 2839
rect 50169 2805 50203 2839
rect 59001 2805 59035 2839
rect 60197 2805 60231 2839
rect 35541 2601 35575 2635
rect 41797 2601 41831 2635
rect 45109 2601 45143 2635
rect 47593 2601 47627 2635
rect 48697 2601 48731 2635
rect 58909 2601 58943 2635
rect 6009 2533 6043 2567
rect 8585 2533 8619 2567
rect 21373 2533 21407 2567
rect 25973 2533 26007 2567
rect 33977 2533 34011 2567
rect 40233 2533 40267 2567
rect 56793 2533 56827 2567
rect 2421 2465 2455 2499
rect 2789 2465 2823 2499
rect 2973 2465 3007 2499
rect 4629 2465 4663 2499
rect 7205 2465 7239 2499
rect 12633 2465 12667 2499
rect 12909 2465 12943 2499
rect 16037 2465 16071 2499
rect 18613 2465 18647 2499
rect 21189 2465 21223 2499
rect 21465 2465 21499 2499
rect 22937 2465 22971 2499
rect 23029 2465 23063 2499
rect 26893 2465 26927 2499
rect 27629 2465 27663 2499
rect 28089 2465 28123 2499
rect 30297 2465 30331 2499
rect 32689 2465 32723 2499
rect 34161 2465 34195 2499
rect 35725 2465 35759 2499
rect 35909 2465 35943 2499
rect 36277 2465 36311 2499
rect 38577 2465 38611 2499
rect 38853 2465 38887 2499
rect 41153 2465 41187 2499
rect 42717 2465 42751 2499
rect 44465 2465 44499 2499
rect 46949 2465 46983 2499
rect 48513 2465 48547 2499
rect 53757 2465 53791 2499
rect 56977 2465 57011 2499
rect 57345 2465 57379 2499
rect 58265 2465 58299 2499
rect 59829 2465 59863 2499
rect 4353 2397 4387 2431
rect 6929 2397 6963 2431
rect 14013 2397 14047 2431
rect 15761 2397 15795 2431
rect 17141 2397 17175 2431
rect 18337 2397 18371 2431
rect 19717 2397 19751 2431
rect 24317 2397 24351 2431
rect 24593 2397 24627 2431
rect 30021 2397 30055 2431
rect 32597 2397 32631 2431
rect 34529 2397 34563 2431
rect 41521 2397 41555 2431
rect 44833 2397 44867 2431
rect 47317 2397 47351 2431
rect 54125 2397 54159 2431
rect 58633 2397 58667 2431
rect 59921 2397 59955 2431
rect 27169 2329 27203 2363
rect 41318 2329 41352 2363
rect 44630 2329 44664 2363
rect 47225 2329 47259 2363
rect 53922 2329 53956 2363
rect 54401 2329 54435 2363
rect 58403 2329 58437 2363
rect 58541 2329 58575 2363
rect 21649 2261 21683 2295
rect 31401 2261 31435 2295
rect 32873 2261 32907 2295
rect 41429 2261 41463 2295
rect 42809 2261 42843 2295
rect 44741 2261 44775 2295
rect 47114 2261 47148 2295
rect 54033 2261 54067 2295
<< metal1 >>
rect 1104 17434 62192 17456
rect 1104 17382 11163 17434
rect 11215 17382 11227 17434
rect 11279 17382 11291 17434
rect 11343 17382 11355 17434
rect 11407 17382 31526 17434
rect 31578 17382 31590 17434
rect 31642 17382 31654 17434
rect 31706 17382 31718 17434
rect 31770 17382 51888 17434
rect 51940 17382 51952 17434
rect 52004 17382 52016 17434
rect 52068 17382 52080 17434
rect 52132 17382 62192 17434
rect 1104 17360 62192 17382
rect 14366 17320 14372 17332
rect 14279 17292 14372 17320
rect 14366 17280 14372 17292
rect 14424 17320 14430 17332
rect 16206 17320 16212 17332
rect 14424 17292 16212 17320
rect 14424 17280 14430 17292
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 19889 17323 19947 17329
rect 19889 17289 19901 17323
rect 19935 17320 19947 17323
rect 20070 17320 20076 17332
rect 19935 17292 20076 17320
rect 19935 17289 19947 17292
rect 19889 17283 19947 17289
rect 20070 17280 20076 17292
rect 20128 17280 20134 17332
rect 25406 17280 25412 17332
rect 25464 17320 25470 17332
rect 25593 17323 25651 17329
rect 25593 17320 25605 17323
rect 25464 17292 25605 17320
rect 25464 17280 25470 17292
rect 25593 17289 25605 17292
rect 25639 17320 25651 17323
rect 27706 17320 27712 17332
rect 25639 17292 27712 17320
rect 25639 17289 25651 17292
rect 25593 17283 25651 17289
rect 27706 17280 27712 17292
rect 27764 17280 27770 17332
rect 40037 17323 40095 17329
rect 40037 17289 40049 17323
rect 40083 17320 40095 17323
rect 40494 17320 40500 17332
rect 40083 17292 40500 17320
rect 40083 17289 40095 17292
rect 40037 17283 40095 17289
rect 40494 17280 40500 17292
rect 40552 17320 40558 17332
rect 41138 17320 41144 17332
rect 40552 17292 41144 17320
rect 40552 17280 40558 17292
rect 41138 17280 41144 17292
rect 41196 17280 41202 17332
rect 45002 17280 45008 17332
rect 45060 17320 45066 17332
rect 45557 17323 45615 17329
rect 45557 17320 45569 17323
rect 45060 17292 45569 17320
rect 45060 17280 45066 17292
rect 45557 17289 45569 17292
rect 45603 17289 45615 17323
rect 45557 17283 45615 17289
rect 11698 17144 11704 17196
rect 11756 17184 11762 17196
rect 12805 17187 12863 17193
rect 12805 17184 12817 17187
rect 11756 17156 12817 17184
rect 11756 17144 11762 17156
rect 12805 17153 12817 17156
rect 12851 17184 12863 17187
rect 16666 17184 16672 17196
rect 12851 17156 16672 17184
rect 12851 17153 12863 17156
rect 12805 17147 12863 17153
rect 16666 17144 16672 17156
rect 16724 17144 16730 17196
rect 25866 17184 25872 17196
rect 22756 17156 25872 17184
rect 13078 17116 13084 17128
rect 13039 17088 13084 17116
rect 13078 17076 13084 17088
rect 13136 17076 13142 17128
rect 16945 17119 17003 17125
rect 16945 17085 16957 17119
rect 16991 17116 17003 17119
rect 17954 17116 17960 17128
rect 16991 17088 17960 17116
rect 16991 17085 17003 17088
rect 16945 17079 17003 17085
rect 17954 17076 17960 17088
rect 18012 17076 18018 17128
rect 18325 17119 18383 17125
rect 18325 17085 18337 17119
rect 18371 17116 18383 17119
rect 18414 17116 18420 17128
rect 18371 17088 18420 17116
rect 18371 17085 18383 17088
rect 18325 17079 18383 17085
rect 18414 17076 18420 17088
rect 18472 17076 18478 17128
rect 18598 17116 18604 17128
rect 18559 17088 18604 17116
rect 18598 17076 18604 17088
rect 18656 17076 18662 17128
rect 22756 17125 22784 17156
rect 25866 17144 25872 17156
rect 25924 17144 25930 17196
rect 37274 17184 37280 17196
rect 35636 17156 37280 17184
rect 22741 17119 22799 17125
rect 22741 17085 22753 17119
rect 22787 17085 22799 17119
rect 24026 17116 24032 17128
rect 23987 17088 24032 17116
rect 22741 17079 22799 17085
rect 24026 17076 24032 17088
rect 24084 17076 24090 17128
rect 24305 17119 24363 17125
rect 24305 17085 24317 17119
rect 24351 17116 24363 17119
rect 24946 17116 24952 17128
rect 24351 17088 24952 17116
rect 24351 17085 24363 17088
rect 24305 17079 24363 17085
rect 24946 17076 24952 17088
rect 25004 17076 25010 17128
rect 28077 17119 28135 17125
rect 28077 17085 28089 17119
rect 28123 17116 28135 17119
rect 29638 17116 29644 17128
rect 28123 17088 29644 17116
rect 28123 17085 28135 17088
rect 28077 17079 28135 17085
rect 29638 17076 29644 17088
rect 29696 17076 29702 17128
rect 33502 17076 33508 17128
rect 33560 17116 33566 17128
rect 35636 17125 35664 17156
rect 37274 17144 37280 17156
rect 37332 17144 37338 17196
rect 37369 17187 37427 17193
rect 37369 17153 37381 17187
rect 37415 17184 37427 17187
rect 38930 17184 38936 17196
rect 37415 17156 38936 17184
rect 37415 17153 37427 17156
rect 37369 17147 37427 17153
rect 38930 17144 38936 17156
rect 38988 17144 38994 17196
rect 34149 17119 34207 17125
rect 34149 17116 34161 17119
rect 33560 17088 34161 17116
rect 33560 17076 33566 17088
rect 34149 17085 34161 17088
rect 34195 17085 34207 17119
rect 34149 17079 34207 17085
rect 35621 17119 35679 17125
rect 35621 17085 35633 17119
rect 35667 17085 35679 17119
rect 35621 17079 35679 17085
rect 37001 17119 37059 17125
rect 37001 17085 37013 17119
rect 37047 17085 37059 17119
rect 37001 17079 37059 17085
rect 15286 17008 15292 17060
rect 15344 17048 15350 17060
rect 16761 17051 16819 17057
rect 16761 17048 16773 17051
rect 15344 17020 16773 17048
rect 15344 17008 15350 17020
rect 16761 17017 16773 17020
rect 16807 17048 16819 17051
rect 17678 17048 17684 17060
rect 16807 17020 17684 17048
rect 16807 17017 16819 17020
rect 16761 17011 16819 17017
rect 17678 17008 17684 17020
rect 17736 17008 17742 17060
rect 22554 17048 22560 17060
rect 22467 17020 22560 17048
rect 22554 17008 22560 17020
rect 22612 17048 22618 17060
rect 22612 17020 24164 17048
rect 22612 17008 22618 17020
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 17037 16983 17095 16989
rect 17037 16980 17049 16983
rect 16632 16952 17049 16980
rect 16632 16940 16638 16952
rect 17037 16949 17049 16952
rect 17083 16949 17095 16983
rect 17037 16943 17095 16949
rect 22186 16940 22192 16992
rect 22244 16980 22250 16992
rect 22833 16983 22891 16989
rect 22833 16980 22845 16983
rect 22244 16952 22845 16980
rect 22244 16940 22250 16952
rect 22833 16949 22845 16952
rect 22879 16949 22891 16983
rect 24136 16980 24164 17020
rect 27246 17008 27252 17060
rect 27304 17048 27310 17060
rect 27893 17051 27951 17057
rect 27893 17048 27905 17051
rect 27304 17020 27905 17048
rect 27304 17008 27310 17020
rect 27893 17017 27905 17020
rect 27939 17048 27951 17051
rect 30190 17048 30196 17060
rect 27939 17020 30196 17048
rect 27939 17017 27951 17020
rect 27893 17011 27951 17017
rect 30190 17008 30196 17020
rect 30248 17008 30254 17060
rect 33965 17051 34023 17057
rect 33965 17017 33977 17051
rect 34011 17048 34023 17051
rect 35437 17051 35495 17057
rect 34011 17020 34928 17048
rect 34011 17017 34023 17020
rect 33965 17011 34023 17017
rect 27264 16980 27292 17008
rect 34900 16992 34928 17020
rect 35437 17017 35449 17051
rect 35483 17017 35495 17051
rect 35986 17048 35992 17060
rect 35947 17020 35992 17048
rect 35437 17011 35495 17017
rect 28166 16980 28172 16992
rect 24136 16952 27292 16980
rect 28127 16952 28172 16980
rect 22833 16943 22891 16949
rect 28166 16940 28172 16952
rect 28224 16940 28230 16992
rect 34238 16980 34244 16992
rect 34199 16952 34244 16980
rect 34238 16940 34244 16952
rect 34296 16940 34302 16992
rect 34882 16940 34888 16992
rect 34940 16980 34946 16992
rect 35452 16980 35480 17011
rect 35986 17008 35992 17020
rect 36044 17008 36050 17060
rect 36814 17048 36820 17060
rect 36775 17020 36820 17048
rect 36814 17008 36820 17020
rect 36872 17008 36878 17060
rect 36832 16980 36860 17008
rect 34940 16952 36860 16980
rect 37016 16980 37044 17079
rect 37826 17076 37832 17128
rect 37884 17116 37890 17128
rect 38473 17119 38531 17125
rect 38473 17116 38485 17119
rect 37884 17088 38485 17116
rect 37884 17076 37890 17088
rect 38473 17085 38485 17088
rect 38519 17085 38531 17119
rect 38746 17116 38752 17128
rect 38707 17088 38752 17116
rect 38473 17079 38531 17085
rect 38746 17076 38752 17088
rect 38804 17076 38810 17128
rect 43990 17116 43996 17128
rect 43951 17088 43996 17116
rect 43990 17076 43996 17088
rect 44048 17076 44054 17128
rect 44266 17116 44272 17128
rect 44227 17088 44272 17116
rect 44266 17076 44272 17088
rect 44324 17076 44330 17128
rect 48409 17119 48467 17125
rect 48409 17085 48421 17119
rect 48455 17116 48467 17119
rect 48866 17116 48872 17128
rect 48455 17088 48872 17116
rect 48455 17085 48467 17088
rect 48409 17079 48467 17085
rect 48866 17076 48872 17088
rect 48924 17076 48930 17128
rect 49881 17119 49939 17125
rect 49881 17085 49893 17119
rect 49927 17116 49939 17119
rect 50798 17116 50804 17128
rect 49927 17088 50804 17116
rect 49927 17085 49939 17088
rect 49881 17079 49939 17085
rect 50798 17076 50804 17088
rect 50856 17076 50862 17128
rect 46198 17008 46204 17060
rect 46256 17048 46262 17060
rect 48225 17051 48283 17057
rect 48225 17048 48237 17051
rect 46256 17020 48237 17048
rect 46256 17008 46262 17020
rect 48225 17017 48237 17020
rect 48271 17048 48283 17051
rect 49697 17051 49755 17057
rect 49697 17048 49709 17051
rect 48271 17020 49709 17048
rect 48271 17017 48283 17020
rect 48225 17011 48283 17017
rect 49697 17017 49709 17020
rect 49743 17017 49755 17051
rect 49697 17011 49755 17017
rect 39206 16980 39212 16992
rect 37016 16952 39212 16980
rect 34940 16940 34946 16952
rect 39206 16940 39212 16952
rect 39264 16940 39270 16992
rect 48498 16980 48504 16992
rect 48459 16952 48504 16980
rect 48498 16940 48504 16952
rect 48556 16940 48562 16992
rect 49970 16980 49976 16992
rect 49931 16952 49976 16980
rect 49970 16940 49976 16952
rect 50028 16940 50034 16992
rect 1104 16890 62192 16912
rect 1104 16838 21344 16890
rect 21396 16838 21408 16890
rect 21460 16838 21472 16890
rect 21524 16838 21536 16890
rect 21588 16838 41707 16890
rect 41759 16838 41771 16890
rect 41823 16838 41835 16890
rect 41887 16838 41899 16890
rect 41951 16838 62192 16890
rect 1104 16816 62192 16838
rect 18049 16779 18107 16785
rect 18049 16776 18061 16779
rect 15488 16748 18061 16776
rect 13449 16711 13507 16717
rect 13449 16677 13461 16711
rect 13495 16708 13507 16711
rect 13814 16708 13820 16720
rect 13495 16680 13820 16708
rect 13495 16677 13507 16680
rect 13449 16671 13507 16677
rect 13814 16668 13820 16680
rect 13872 16708 13878 16720
rect 14274 16708 14280 16720
rect 13872 16680 14280 16708
rect 13872 16668 13878 16680
rect 14274 16668 14280 16680
rect 14332 16668 14338 16720
rect 15286 16708 15292 16720
rect 15247 16680 15292 16708
rect 15286 16668 15292 16680
rect 15344 16668 15350 16720
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 11793 16643 11851 16649
rect 11793 16640 11805 16643
rect 11756 16612 11805 16640
rect 11756 16600 11762 16612
rect 11793 16609 11805 16612
rect 11839 16609 11851 16643
rect 11793 16603 11851 16609
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16640 12127 16643
rect 12526 16640 12532 16652
rect 12115 16612 12532 16640
rect 12115 16609 12127 16612
rect 12069 16603 12127 16609
rect 12526 16600 12532 16612
rect 12584 16600 12590 16652
rect 15488 16649 15516 16748
rect 18049 16745 18061 16748
rect 18095 16776 18107 16779
rect 18138 16776 18144 16788
rect 18095 16748 18144 16776
rect 18095 16745 18107 16748
rect 18049 16739 18107 16745
rect 18138 16736 18144 16748
rect 18196 16736 18202 16788
rect 23934 16736 23940 16788
rect 23992 16776 23998 16788
rect 24121 16779 24179 16785
rect 24121 16776 24133 16779
rect 23992 16748 24133 16776
rect 23992 16736 23998 16748
rect 24121 16745 24133 16748
rect 24167 16745 24179 16779
rect 24121 16739 24179 16745
rect 33502 16736 33508 16788
rect 33560 16776 33566 16788
rect 33781 16779 33839 16785
rect 33781 16776 33793 16779
rect 33560 16748 33793 16776
rect 33560 16736 33566 16748
rect 33781 16745 33793 16748
rect 33827 16745 33839 16779
rect 33781 16739 33839 16745
rect 36814 16736 36820 16788
rect 36872 16776 36878 16788
rect 39206 16776 39212 16788
rect 36872 16748 38792 16776
rect 39167 16748 39212 16776
rect 36872 16736 36878 16748
rect 17678 16668 17684 16720
rect 17736 16708 17742 16720
rect 19153 16711 19211 16717
rect 19153 16708 19165 16711
rect 17736 16680 19165 16708
rect 17736 16668 17742 16680
rect 19153 16677 19165 16680
rect 19199 16677 19211 16711
rect 19153 16671 19211 16677
rect 21361 16711 21419 16717
rect 21361 16677 21373 16711
rect 21407 16708 21419 16711
rect 22554 16708 22560 16720
rect 21407 16680 22560 16708
rect 21407 16677 21419 16680
rect 21361 16671 21419 16677
rect 22554 16668 22560 16680
rect 22612 16668 22618 16720
rect 15473 16643 15531 16649
rect 15473 16609 15485 16643
rect 15519 16609 15531 16643
rect 16666 16640 16672 16652
rect 16627 16612 16672 16640
rect 15473 16603 15531 16609
rect 16666 16600 16672 16612
rect 16724 16600 16730 16652
rect 16942 16640 16948 16652
rect 16903 16612 16948 16640
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 19337 16643 19395 16649
rect 19337 16609 19349 16643
rect 19383 16640 19395 16643
rect 20070 16640 20076 16652
rect 19383 16612 20076 16640
rect 19383 16609 19395 16612
rect 19337 16603 19395 16609
rect 20070 16600 20076 16612
rect 20128 16600 20134 16652
rect 21545 16643 21603 16649
rect 21545 16609 21557 16643
rect 21591 16640 21603 16643
rect 23952 16640 23980 16736
rect 29365 16711 29423 16717
rect 29365 16677 29377 16711
rect 29411 16708 29423 16711
rect 29638 16708 29644 16720
rect 29411 16680 29644 16708
rect 29411 16677 29423 16680
rect 29365 16671 29423 16677
rect 29638 16668 29644 16680
rect 29696 16668 29702 16720
rect 30190 16708 30196 16720
rect 30151 16680 30196 16708
rect 30190 16668 30196 16680
rect 30248 16668 30254 16720
rect 38764 16708 38792 16748
rect 39206 16736 39212 16748
rect 39264 16736 39270 16788
rect 46934 16736 46940 16788
rect 46992 16776 46998 16788
rect 47213 16779 47271 16785
rect 47213 16776 47225 16779
rect 46992 16748 47225 16776
rect 46992 16736 46998 16748
rect 47213 16745 47225 16748
rect 47259 16745 47271 16779
rect 50798 16776 50804 16788
rect 50759 16748 50804 16776
rect 47213 16739 47271 16745
rect 50798 16736 50804 16748
rect 50856 16736 50862 16788
rect 40313 16711 40371 16717
rect 40313 16708 40325 16711
rect 38764 16680 40325 16708
rect 40313 16677 40325 16680
rect 40359 16677 40371 16711
rect 40313 16671 40371 16677
rect 56965 16711 57023 16717
rect 56965 16677 56977 16711
rect 57011 16708 57023 16711
rect 57011 16680 57100 16708
rect 57011 16677 57023 16680
rect 56965 16671 57023 16677
rect 21591 16612 23980 16640
rect 27709 16643 27767 16649
rect 21591 16609 21603 16612
rect 21545 16603 21603 16609
rect 27709 16609 27721 16643
rect 27755 16640 27767 16643
rect 29270 16640 29276 16652
rect 27755 16612 29276 16640
rect 27755 16609 27767 16612
rect 27709 16603 27767 16609
rect 29270 16600 29276 16612
rect 29328 16600 29334 16652
rect 30377 16643 30435 16649
rect 30377 16609 30389 16643
rect 30423 16640 30435 16643
rect 31386 16640 31392 16652
rect 30423 16612 31392 16640
rect 30423 16609 30435 16612
rect 30377 16603 30435 16609
rect 31386 16600 31392 16612
rect 31444 16600 31450 16652
rect 32677 16643 32735 16649
rect 32677 16609 32689 16643
rect 32723 16640 32735 16643
rect 34790 16640 34796 16652
rect 32723 16612 34796 16640
rect 32723 16609 32735 16612
rect 32677 16603 32735 16609
rect 34790 16600 34796 16612
rect 34848 16600 34854 16652
rect 35158 16640 35164 16652
rect 35119 16612 35164 16640
rect 35158 16600 35164 16612
rect 35216 16600 35222 16652
rect 37826 16640 37832 16652
rect 37787 16612 37832 16640
rect 37826 16600 37832 16612
rect 37884 16600 37890 16652
rect 38105 16643 38163 16649
rect 38105 16609 38117 16643
rect 38151 16640 38163 16643
rect 39206 16640 39212 16652
rect 38151 16612 39212 16640
rect 38151 16609 38163 16612
rect 38105 16603 38163 16609
rect 39206 16600 39212 16612
rect 39264 16600 39270 16652
rect 40494 16640 40500 16652
rect 40455 16612 40500 16640
rect 40494 16600 40500 16612
rect 40552 16600 40558 16652
rect 42886 16600 42892 16652
rect 42944 16640 42950 16652
rect 43349 16643 43407 16649
rect 43349 16640 43361 16643
rect 42944 16612 43361 16640
rect 42944 16600 42950 16612
rect 43349 16609 43361 16612
rect 43395 16640 43407 16643
rect 43990 16640 43996 16652
rect 43395 16612 43996 16640
rect 43395 16609 43407 16612
rect 43349 16603 43407 16609
rect 43990 16600 43996 16612
rect 44048 16600 44054 16652
rect 45833 16643 45891 16649
rect 45833 16609 45845 16643
rect 45879 16640 45891 16643
rect 45922 16640 45928 16652
rect 45879 16612 45928 16640
rect 45879 16609 45891 16612
rect 45833 16603 45891 16609
rect 45922 16600 45928 16612
rect 45980 16640 45986 16652
rect 48038 16640 48044 16652
rect 45980 16612 48044 16640
rect 45980 16600 45986 16612
rect 48038 16600 48044 16612
rect 48096 16640 48102 16652
rect 49421 16643 49479 16649
rect 49421 16640 49433 16643
rect 48096 16612 49433 16640
rect 48096 16600 48102 16612
rect 49421 16609 49433 16612
rect 49467 16609 49479 16643
rect 55306 16640 55312 16652
rect 55267 16612 55312 16640
rect 49421 16603 49479 16609
rect 55306 16600 55312 16612
rect 55364 16600 55370 16652
rect 55582 16640 55588 16652
rect 55543 16612 55588 16640
rect 55582 16600 55588 16612
rect 55640 16600 55646 16652
rect 57072 16584 57100 16680
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16572 15899 16575
rect 16482 16572 16488 16584
rect 15887 16544 16488 16572
rect 15887 16541 15899 16544
rect 15841 16535 15899 16541
rect 16482 16532 16488 16544
rect 16540 16532 16546 16584
rect 18414 16532 18420 16584
rect 18472 16572 18478 16584
rect 22738 16572 22744 16584
rect 18472 16544 22744 16572
rect 18472 16532 18478 16544
rect 22738 16532 22744 16544
rect 22796 16532 22802 16584
rect 23014 16572 23020 16584
rect 22975 16544 23020 16572
rect 23014 16532 23020 16544
rect 23072 16532 23078 16584
rect 27982 16572 27988 16584
rect 27943 16544 27988 16572
rect 27982 16532 27988 16544
rect 28040 16532 28046 16584
rect 32401 16575 32459 16581
rect 32401 16541 32413 16575
rect 32447 16572 32459 16575
rect 32858 16572 32864 16584
rect 32447 16544 32864 16572
rect 32447 16541 32459 16544
rect 32401 16535 32459 16541
rect 32858 16532 32864 16544
rect 32916 16572 32922 16584
rect 34885 16575 34943 16581
rect 34885 16572 34897 16575
rect 32916 16544 34897 16572
rect 32916 16532 32922 16544
rect 34885 16541 34897 16544
rect 34931 16572 34943 16575
rect 35250 16572 35256 16584
rect 34931 16544 35256 16572
rect 34931 16541 34943 16544
rect 34885 16535 34943 16541
rect 35250 16532 35256 16544
rect 35308 16532 35314 16584
rect 35526 16532 35532 16584
rect 35584 16572 35590 16584
rect 36265 16575 36323 16581
rect 36265 16572 36277 16575
rect 35584 16544 36277 16572
rect 35584 16532 35590 16544
rect 36265 16541 36277 16544
rect 36311 16541 36323 16575
rect 36265 16535 36323 16541
rect 43625 16575 43683 16581
rect 43625 16541 43637 16575
rect 43671 16572 43683 16575
rect 43714 16572 43720 16584
rect 43671 16544 43720 16572
rect 43671 16541 43683 16544
rect 43625 16535 43683 16541
rect 43714 16532 43720 16544
rect 43772 16532 43778 16584
rect 46106 16572 46112 16584
rect 46067 16544 46112 16572
rect 46106 16532 46112 16544
rect 46164 16532 46170 16584
rect 49694 16572 49700 16584
rect 49655 16544 49700 16572
rect 49694 16532 49700 16544
rect 49752 16532 49758 16584
rect 57054 16532 57060 16584
rect 57112 16572 57118 16584
rect 58434 16572 58440 16584
rect 57112 16544 58440 16572
rect 57112 16532 57118 16544
rect 58434 16532 58440 16544
rect 58492 16532 58498 16584
rect 18230 16396 18236 16448
rect 18288 16436 18294 16448
rect 19429 16439 19487 16445
rect 19429 16436 19441 16439
rect 18288 16408 19441 16436
rect 18288 16396 18294 16408
rect 19429 16405 19441 16408
rect 19475 16405 19487 16439
rect 19429 16399 19487 16405
rect 21637 16439 21695 16445
rect 21637 16405 21649 16439
rect 21683 16436 21695 16439
rect 22922 16436 22928 16448
rect 21683 16408 22928 16436
rect 21683 16405 21695 16408
rect 21637 16399 21695 16405
rect 22922 16396 22928 16408
rect 22980 16396 22986 16448
rect 28718 16396 28724 16448
rect 28776 16436 28782 16448
rect 30469 16439 30527 16445
rect 30469 16436 30481 16439
rect 28776 16408 30481 16436
rect 28776 16396 28782 16408
rect 30469 16405 30481 16408
rect 30515 16405 30527 16439
rect 40586 16436 40592 16448
rect 40547 16408 40592 16436
rect 30469 16399 30527 16405
rect 40586 16396 40592 16408
rect 40644 16396 40650 16448
rect 43070 16396 43076 16448
rect 43128 16436 43134 16448
rect 44729 16439 44787 16445
rect 44729 16436 44741 16439
rect 43128 16408 44741 16436
rect 43128 16396 43134 16408
rect 44729 16405 44741 16408
rect 44775 16405 44787 16439
rect 44729 16399 44787 16405
rect 1104 16346 62192 16368
rect 1104 16294 11163 16346
rect 11215 16294 11227 16346
rect 11279 16294 11291 16346
rect 11343 16294 11355 16346
rect 11407 16294 31526 16346
rect 31578 16294 31590 16346
rect 31642 16294 31654 16346
rect 31706 16294 31718 16346
rect 31770 16294 51888 16346
rect 51940 16294 51952 16346
rect 52004 16294 52016 16346
rect 52068 16294 52080 16346
rect 52132 16294 62192 16346
rect 1104 16272 62192 16294
rect 13078 16232 13084 16244
rect 13039 16204 13084 16232
rect 13078 16192 13084 16204
rect 13136 16192 13142 16244
rect 18509 16235 18567 16241
rect 18509 16201 18521 16235
rect 18555 16232 18567 16235
rect 18598 16232 18604 16244
rect 18555 16204 18604 16232
rect 18555 16201 18567 16204
rect 18509 16195 18567 16201
rect 18598 16192 18604 16204
rect 18656 16192 18662 16244
rect 22005 16235 22063 16241
rect 22005 16201 22017 16235
rect 22051 16232 22063 16235
rect 23658 16232 23664 16244
rect 22051 16204 23664 16232
rect 22051 16201 22063 16204
rect 22005 16195 22063 16201
rect 23658 16192 23664 16204
rect 23716 16232 23722 16244
rect 25225 16235 25283 16241
rect 23716 16204 25176 16232
rect 23716 16192 23722 16204
rect 12621 16167 12679 16173
rect 12621 16133 12633 16167
rect 12667 16164 12679 16167
rect 16209 16167 16267 16173
rect 16209 16164 16221 16167
rect 12667 16136 16221 16164
rect 12667 16133 12679 16136
rect 12621 16127 12679 16133
rect 16209 16133 16221 16136
rect 16255 16164 16267 16167
rect 16298 16164 16304 16176
rect 16255 16136 16304 16164
rect 16255 16133 16267 16136
rect 16209 16127 16267 16133
rect 12158 15988 12164 16040
rect 12216 16028 12222 16040
rect 12636 16028 12664 16127
rect 16298 16124 16304 16136
rect 16356 16164 16362 16176
rect 18049 16167 18107 16173
rect 18049 16164 18061 16167
rect 16356 16136 18061 16164
rect 16356 16124 16362 16136
rect 18049 16133 18061 16136
rect 18095 16133 18107 16167
rect 25148 16164 25176 16204
rect 25225 16201 25237 16235
rect 25271 16232 25283 16235
rect 25866 16232 25872 16244
rect 25271 16204 25872 16232
rect 25271 16201 25283 16204
rect 25225 16195 25283 16201
rect 25866 16192 25872 16204
rect 25924 16192 25930 16244
rect 30837 16235 30895 16241
rect 30837 16201 30849 16235
rect 30883 16232 30895 16235
rect 31386 16232 31392 16244
rect 30883 16204 31392 16232
rect 30883 16201 30895 16204
rect 30837 16195 30895 16201
rect 31386 16192 31392 16204
rect 31444 16192 31450 16244
rect 33873 16235 33931 16241
rect 33873 16201 33885 16235
rect 33919 16232 33931 16235
rect 34882 16232 34888 16244
rect 33919 16204 34888 16232
rect 33919 16201 33931 16204
rect 33873 16195 33931 16201
rect 34882 16192 34888 16204
rect 34940 16192 34946 16244
rect 37366 16192 37372 16244
rect 37424 16232 37430 16244
rect 37645 16235 37703 16241
rect 37645 16232 37657 16235
rect 37424 16204 37657 16232
rect 37424 16192 37430 16204
rect 37645 16201 37657 16204
rect 37691 16201 37703 16235
rect 39206 16232 39212 16244
rect 39167 16204 39212 16232
rect 37645 16195 37703 16201
rect 39206 16192 39212 16204
rect 39264 16192 39270 16244
rect 44266 16192 44272 16244
rect 44324 16232 44330 16244
rect 44729 16235 44787 16241
rect 44729 16232 44741 16235
rect 44324 16204 44741 16232
rect 44324 16192 44330 16204
rect 44729 16201 44741 16204
rect 44775 16201 44787 16235
rect 44729 16195 44787 16201
rect 48958 16192 48964 16244
rect 49016 16232 49022 16244
rect 49421 16235 49479 16241
rect 49421 16232 49433 16235
rect 49016 16204 49433 16232
rect 49016 16192 49022 16204
rect 49421 16201 49433 16204
rect 49467 16201 49479 16235
rect 49421 16195 49479 16201
rect 27249 16167 27307 16173
rect 27249 16164 27261 16167
rect 25148 16136 27261 16164
rect 18049 16127 18107 16133
rect 27249 16133 27261 16136
rect 27295 16164 27307 16167
rect 27890 16164 27896 16176
rect 27295 16136 27896 16164
rect 27295 16133 27307 16136
rect 27249 16127 27307 16133
rect 27890 16124 27896 16136
rect 27948 16124 27954 16176
rect 41969 16167 42027 16173
rect 41969 16133 41981 16167
rect 42015 16164 42027 16167
rect 42015 16136 42932 16164
rect 42015 16133 42027 16136
rect 41969 16127 42027 16133
rect 15470 16056 15476 16108
rect 15528 16096 15534 16108
rect 22741 16099 22799 16105
rect 15528 16068 22692 16096
rect 15528 16056 15534 16068
rect 12216 16000 12664 16028
rect 12216 15988 12222 16000
rect 12710 15988 12716 16040
rect 12768 16028 12774 16040
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 12768 16000 12909 16028
rect 12768 15988 12774 16000
rect 12897 15997 12909 16000
rect 12943 15997 12955 16031
rect 14366 16028 14372 16040
rect 14327 16000 14372 16028
rect 12897 15991 12955 15997
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 15194 15988 15200 16040
rect 15252 16028 15258 16040
rect 16485 16031 16543 16037
rect 16485 16028 16497 16031
rect 15252 16000 16497 16028
rect 15252 15988 15258 16000
rect 16485 15997 16497 16000
rect 16531 15997 16543 16031
rect 18230 16028 18236 16040
rect 18191 16000 18236 16028
rect 16485 15991 16543 15997
rect 18230 15988 18236 16000
rect 18288 15988 18294 16040
rect 18322 15988 18328 16040
rect 18380 16028 18386 16040
rect 20622 16028 20628 16040
rect 18380 16000 18425 16028
rect 20583 16000 20628 16028
rect 18380 15988 18386 16000
rect 20622 15988 20628 16000
rect 20680 15988 20686 16040
rect 20717 16031 20775 16037
rect 20717 15997 20729 16031
rect 20763 15997 20775 16031
rect 22278 16028 22284 16040
rect 22239 16000 22284 16028
rect 20717 15991 20775 15997
rect 2774 15920 2780 15972
rect 2832 15960 2838 15972
rect 12342 15960 12348 15972
rect 2832 15932 12348 15960
rect 2832 15920 2838 15932
rect 12342 15920 12348 15932
rect 12400 15920 12406 15972
rect 12805 15963 12863 15969
rect 12805 15929 12817 15963
rect 12851 15929 12863 15963
rect 12805 15923 12863 15929
rect 14185 15963 14243 15969
rect 14185 15929 14197 15963
rect 14231 15960 14243 15963
rect 15286 15960 15292 15972
rect 14231 15932 15292 15960
rect 14231 15929 14243 15932
rect 14185 15923 14243 15929
rect 934 15852 940 15904
rect 992 15892 998 15904
rect 10134 15892 10140 15904
rect 992 15864 10140 15892
rect 992 15852 998 15864
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 12820 15892 12848 15923
rect 15286 15920 15292 15932
rect 15344 15920 15350 15972
rect 16393 15963 16451 15969
rect 16393 15929 16405 15963
rect 16439 15960 16451 15963
rect 16574 15960 16580 15972
rect 16439 15932 16580 15960
rect 16439 15929 16451 15932
rect 16393 15923 16451 15929
rect 16574 15920 16580 15932
rect 16632 15920 16638 15972
rect 16945 15963 17003 15969
rect 16945 15929 16957 15963
rect 16991 15960 17003 15963
rect 17218 15960 17224 15972
rect 16991 15932 17224 15960
rect 16991 15929 17003 15932
rect 16945 15923 17003 15929
rect 17218 15920 17224 15932
rect 17276 15920 17282 15972
rect 19518 15920 19524 15972
rect 19576 15960 19582 15972
rect 20732 15960 20760 15991
rect 22278 15988 22284 16000
rect 22336 15988 22342 16040
rect 21174 15960 21180 15972
rect 19576 15932 20760 15960
rect 21135 15932 21180 15960
rect 19576 15920 19582 15932
rect 21174 15920 21180 15932
rect 21232 15920 21238 15972
rect 22186 15960 22192 15972
rect 22147 15932 22192 15960
rect 22186 15920 22192 15932
rect 22244 15920 22250 15972
rect 14461 15895 14519 15901
rect 14461 15892 14473 15895
rect 12820 15864 14473 15892
rect 14461 15861 14473 15864
rect 14507 15861 14519 15895
rect 22664 15892 22692 16068
rect 22741 16065 22753 16099
rect 22787 16096 22799 16099
rect 23937 16099 23995 16105
rect 23937 16096 23949 16099
rect 22787 16068 23949 16096
rect 22787 16065 22799 16068
rect 22741 16059 22799 16065
rect 23937 16065 23949 16068
rect 23983 16065 23995 16099
rect 27982 16096 27988 16108
rect 27943 16068 27988 16096
rect 23937 16059 23995 16065
rect 27982 16056 27988 16068
rect 28040 16056 28046 16108
rect 35250 16056 35256 16108
rect 35308 16096 35314 16108
rect 36265 16099 36323 16105
rect 36265 16096 36277 16099
rect 35308 16068 36277 16096
rect 35308 16056 35314 16068
rect 36265 16065 36277 16068
rect 36311 16096 36323 16099
rect 37826 16096 37832 16108
rect 36311 16068 37832 16096
rect 36311 16065 36323 16068
rect 36265 16059 36323 16065
rect 37826 16056 37832 16068
rect 37884 16056 37890 16108
rect 42904 16096 42932 16136
rect 42904 16068 44772 16096
rect 22830 15988 22836 16040
rect 22888 16028 22894 16040
rect 23661 16031 23719 16037
rect 23661 16028 23673 16031
rect 22888 16000 23673 16028
rect 22888 15988 22894 16000
rect 23661 15997 23673 16000
rect 23707 16028 23719 16031
rect 24026 16028 24032 16040
rect 23707 16000 24032 16028
rect 23707 15997 23719 16000
rect 23661 15991 23719 15997
rect 24026 15988 24032 16000
rect 24084 15988 24090 16040
rect 27525 16031 27583 16037
rect 27525 16028 27537 16031
rect 27356 16000 27537 16028
rect 24854 15920 24860 15972
rect 24912 15960 24918 15972
rect 27356 15960 27384 16000
rect 27525 15997 27537 16000
rect 27571 15997 27583 16031
rect 29270 16028 29276 16040
rect 29231 16000 29276 16028
rect 27525 15991 27583 15997
rect 29270 15988 29276 16000
rect 29328 15988 29334 16040
rect 29546 16028 29552 16040
rect 29507 16000 29552 16028
rect 29546 15988 29552 16000
rect 29604 15988 29610 16040
rect 33689 16031 33747 16037
rect 33689 15997 33701 16031
rect 33735 16028 33747 16031
rect 33870 16028 33876 16040
rect 33735 16000 33876 16028
rect 33735 15997 33747 16000
rect 33689 15991 33747 15997
rect 33870 15988 33876 16000
rect 33928 15988 33934 16040
rect 34882 16028 34888 16040
rect 34843 16000 34888 16028
rect 34882 15988 34888 16000
rect 34940 15988 34946 16040
rect 35069 16031 35127 16037
rect 35069 15997 35081 16031
rect 35115 16028 35127 16031
rect 35526 16028 35532 16040
rect 35115 16000 35532 16028
rect 35115 15997 35127 16000
rect 35069 15991 35127 15997
rect 35526 15988 35532 16000
rect 35584 15988 35590 16040
rect 36538 16028 36544 16040
rect 36499 16000 36544 16028
rect 36538 15988 36544 16000
rect 36596 15988 36602 16040
rect 38378 15988 38384 16040
rect 38436 16028 38442 16040
rect 38749 16031 38807 16037
rect 38749 16028 38761 16031
rect 38436 16000 38761 16028
rect 38436 15988 38442 16000
rect 38749 15997 38761 16000
rect 38795 15997 38807 16031
rect 38930 16028 38936 16040
rect 38891 16000 38936 16028
rect 38749 15991 38807 15997
rect 38930 15988 38936 16000
rect 38988 15988 38994 16040
rect 39025 16031 39083 16037
rect 39025 15997 39037 16031
rect 39071 15997 39083 16031
rect 39025 15991 39083 15997
rect 41785 16031 41843 16037
rect 41785 15997 41797 16031
rect 41831 16028 41843 16031
rect 42058 16028 42064 16040
rect 41831 16000 42064 16028
rect 41831 15997 41843 16000
rect 41785 15991 41843 15997
rect 24912 15932 27384 15960
rect 27433 15963 27491 15969
rect 24912 15920 24918 15932
rect 27433 15929 27445 15963
rect 27479 15960 27491 15963
rect 28166 15960 28172 15972
rect 27479 15932 28172 15960
rect 27479 15929 27491 15932
rect 27433 15923 27491 15929
rect 28166 15920 28172 15932
rect 28224 15920 28230 15972
rect 35342 15920 35348 15972
rect 35400 15960 35406 15972
rect 35437 15963 35495 15969
rect 35437 15960 35449 15963
rect 35400 15932 35449 15960
rect 35400 15920 35406 15932
rect 35437 15929 35449 15932
rect 35483 15929 35495 15963
rect 35437 15923 35495 15929
rect 38194 15920 38200 15972
rect 38252 15960 38258 15972
rect 39040 15960 39068 15991
rect 42058 15988 42064 16000
rect 42116 15988 42122 16040
rect 42904 16037 42932 16068
rect 44744 16040 44772 16068
rect 46658 16056 46664 16108
rect 46716 16096 46722 16108
rect 62298 16096 62304 16108
rect 46716 16068 62304 16096
rect 46716 16056 46722 16068
rect 62298 16056 62304 16068
rect 62356 16056 62362 16108
rect 42889 16031 42947 16037
rect 42889 15997 42901 16031
rect 42935 15997 42947 16031
rect 43070 16028 43076 16040
rect 43031 16000 43076 16028
rect 42889 15991 42947 15997
rect 43070 15988 43076 16000
rect 43128 15988 43134 16040
rect 44082 15988 44088 16040
rect 44140 16028 44146 16040
rect 44269 16031 44327 16037
rect 44269 16028 44281 16031
rect 44140 16000 44281 16028
rect 44140 15988 44146 16000
rect 44269 15997 44281 16000
rect 44315 15997 44327 16031
rect 44542 16028 44548 16040
rect 44503 16000 44548 16028
rect 44269 15991 44327 15997
rect 44542 15988 44548 16000
rect 44600 15988 44606 16040
rect 44726 15988 44732 16040
rect 44784 16028 44790 16040
rect 46109 16031 46167 16037
rect 46109 16028 46121 16031
rect 44784 16000 46121 16028
rect 44784 15988 44790 16000
rect 46109 15997 46121 16000
rect 46155 16028 46167 16031
rect 46198 16028 46204 16040
rect 46155 16000 46204 16028
rect 46155 15997 46167 16000
rect 46109 15991 46167 15997
rect 46198 15988 46204 16000
rect 46256 15988 46262 16040
rect 46293 16031 46351 16037
rect 46293 15997 46305 16031
rect 46339 16028 46351 16031
rect 46934 16028 46940 16040
rect 46339 16000 46940 16028
rect 46339 15997 46351 16000
rect 46293 15991 46351 15997
rect 46934 15988 46940 16000
rect 46992 15988 46998 16040
rect 48038 16028 48044 16040
rect 47999 16000 48044 16028
rect 48038 15988 48044 16000
rect 48096 15988 48102 16040
rect 48314 16028 48320 16040
rect 48275 16000 48320 16028
rect 48314 15988 48320 16000
rect 48372 15988 48378 16040
rect 55769 16031 55827 16037
rect 55769 15997 55781 16031
rect 55815 16028 55827 16031
rect 57054 16028 57060 16040
rect 55815 16000 57060 16028
rect 55815 15997 55827 16000
rect 55769 15991 55827 15997
rect 57054 15988 57060 16000
rect 57112 15988 57118 16040
rect 38252 15932 39068 15960
rect 43441 15963 43499 15969
rect 38252 15920 38258 15932
rect 43441 15929 43453 15963
rect 43487 15960 43499 15963
rect 43622 15960 43628 15972
rect 43487 15932 43628 15960
rect 43487 15929 43499 15932
rect 43441 15923 43499 15929
rect 43622 15920 43628 15932
rect 43680 15920 43686 15972
rect 44450 15960 44456 15972
rect 44411 15932 44456 15960
rect 44450 15920 44456 15932
rect 44508 15920 44514 15972
rect 55122 15920 55128 15972
rect 55180 15960 55186 15972
rect 55585 15963 55643 15969
rect 55585 15960 55597 15963
rect 55180 15932 55597 15960
rect 55180 15920 55186 15932
rect 55585 15929 55597 15932
rect 55631 15929 55643 15963
rect 55585 15923 55643 15929
rect 27062 15892 27068 15904
rect 22664 15864 27068 15892
rect 14461 15855 14519 15861
rect 27062 15852 27068 15864
rect 27120 15852 27126 15904
rect 45186 15852 45192 15904
rect 45244 15892 45250 15904
rect 46385 15895 46443 15901
rect 46385 15892 46397 15895
rect 45244 15864 46397 15892
rect 45244 15852 45250 15864
rect 46385 15861 46397 15864
rect 46431 15861 46443 15895
rect 55858 15892 55864 15904
rect 55819 15864 55864 15892
rect 46385 15855 46443 15861
rect 55858 15852 55864 15864
rect 55916 15852 55922 15904
rect 1104 15802 62192 15824
rect 1104 15750 21344 15802
rect 21396 15750 21408 15802
rect 21460 15750 21472 15802
rect 21524 15750 21536 15802
rect 21588 15750 41707 15802
rect 41759 15750 41771 15802
rect 41823 15750 41835 15802
rect 41887 15750 41899 15802
rect 41951 15750 62192 15802
rect 1104 15728 62192 15750
rect 12342 15648 12348 15700
rect 12400 15688 12406 15700
rect 22097 15691 22155 15697
rect 22097 15688 22109 15691
rect 12400 15660 22109 15688
rect 12400 15648 12406 15660
rect 22097 15657 22109 15660
rect 22143 15657 22155 15691
rect 22097 15651 22155 15657
rect 27062 15648 27068 15700
rect 27120 15688 27126 15700
rect 33870 15688 33876 15700
rect 27120 15660 33876 15688
rect 27120 15648 27126 15660
rect 33870 15648 33876 15660
rect 33928 15648 33934 15700
rect 36078 15648 36084 15700
rect 36136 15688 36142 15700
rect 38378 15688 38384 15700
rect 36136 15660 38384 15688
rect 36136 15648 36142 15660
rect 38378 15648 38384 15660
rect 38436 15648 38442 15700
rect 48498 15688 48504 15700
rect 47504 15660 48504 15688
rect 4706 15580 4712 15632
rect 4764 15620 4770 15632
rect 7469 15623 7527 15629
rect 4764 15592 5764 15620
rect 4764 15580 4770 15592
rect 5736 15561 5764 15592
rect 7469 15589 7481 15623
rect 7515 15620 7527 15623
rect 8110 15620 8116 15632
rect 7515 15592 8116 15620
rect 7515 15589 7527 15592
rect 7469 15583 7527 15589
rect 5537 15555 5595 15561
rect 5537 15521 5549 15555
rect 5583 15521 5595 15555
rect 5537 15515 5595 15521
rect 5721 15555 5779 15561
rect 5721 15521 5733 15555
rect 5767 15552 5779 15555
rect 5994 15552 6000 15564
rect 5767 15524 6000 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 5442 15444 5448 15496
rect 5500 15484 5506 15496
rect 5552 15484 5580 15515
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 7484 15484 7512 15583
rect 8110 15580 8116 15592
rect 8168 15580 8174 15632
rect 12253 15623 12311 15629
rect 12253 15589 12265 15623
rect 12299 15620 12311 15623
rect 14185 15623 14243 15629
rect 14185 15620 14197 15623
rect 12299 15592 14197 15620
rect 12299 15589 12311 15592
rect 12253 15583 12311 15589
rect 14185 15589 14197 15592
rect 14231 15589 14243 15623
rect 14185 15583 14243 15589
rect 17954 15580 17960 15632
rect 18012 15620 18018 15632
rect 18601 15623 18659 15629
rect 18601 15620 18613 15623
rect 18012 15592 18613 15620
rect 18012 15580 18018 15592
rect 18601 15589 18613 15592
rect 18647 15620 18659 15623
rect 22002 15620 22008 15632
rect 18647 15592 22008 15620
rect 18647 15589 18659 15592
rect 18601 15583 18659 15589
rect 22002 15580 22008 15592
rect 22060 15580 22066 15632
rect 22189 15623 22247 15629
rect 22189 15589 22201 15623
rect 22235 15620 22247 15623
rect 22278 15620 22284 15632
rect 22235 15592 22284 15620
rect 22235 15589 22247 15592
rect 22189 15583 22247 15589
rect 22278 15580 22284 15592
rect 22336 15580 22342 15632
rect 24946 15620 24952 15632
rect 24907 15592 24952 15620
rect 24946 15580 24952 15592
rect 25004 15580 25010 15632
rect 28718 15620 28724 15632
rect 28679 15592 28724 15620
rect 28718 15580 28724 15592
rect 28776 15580 28782 15632
rect 29273 15623 29331 15629
rect 29273 15589 29285 15623
rect 29319 15620 29331 15623
rect 29546 15620 29552 15632
rect 29319 15592 29552 15620
rect 29319 15589 29331 15592
rect 29273 15583 29331 15589
rect 29546 15580 29552 15592
rect 29604 15580 29610 15632
rect 35986 15580 35992 15632
rect 36044 15620 36050 15632
rect 36265 15623 36323 15629
rect 36265 15620 36277 15623
rect 36044 15592 36277 15620
rect 36044 15580 36050 15592
rect 36265 15589 36277 15592
rect 36311 15589 36323 15623
rect 36265 15583 36323 15589
rect 38473 15623 38531 15629
rect 38473 15589 38485 15623
rect 38519 15620 38531 15623
rect 40586 15620 40592 15632
rect 38519 15592 40592 15620
rect 38519 15589 38531 15592
rect 38473 15583 38531 15589
rect 40586 15580 40592 15592
rect 40644 15580 40650 15632
rect 43622 15620 43628 15632
rect 43583 15592 43628 15620
rect 43622 15580 43628 15592
rect 43680 15580 43686 15632
rect 45186 15620 45192 15632
rect 45147 15592 45192 15620
rect 45186 15580 45192 15592
rect 45244 15580 45250 15632
rect 45741 15623 45799 15629
rect 45741 15589 45753 15623
rect 45787 15620 45799 15623
rect 46106 15620 46112 15632
rect 45787 15592 46112 15620
rect 45787 15589 45799 15592
rect 45741 15583 45799 15589
rect 46106 15580 46112 15592
rect 46164 15580 46170 15632
rect 47504 15629 47532 15660
rect 48498 15648 48504 15660
rect 48556 15648 48562 15700
rect 49970 15688 49976 15700
rect 49160 15660 49976 15688
rect 47489 15623 47547 15629
rect 47489 15589 47501 15623
rect 47535 15589 47547 15623
rect 47489 15583 47547 15589
rect 48041 15623 48099 15629
rect 48041 15589 48053 15623
rect 48087 15620 48099 15623
rect 48314 15620 48320 15632
rect 48087 15592 48320 15620
rect 48087 15589 48099 15592
rect 48041 15583 48099 15589
rect 48314 15580 48320 15592
rect 48372 15580 48378 15632
rect 49160 15629 49188 15660
rect 49970 15648 49976 15660
rect 50028 15648 50034 15700
rect 49145 15623 49203 15629
rect 49145 15589 49157 15623
rect 49191 15589 49203 15623
rect 49694 15620 49700 15632
rect 49655 15592 49700 15620
rect 49145 15583 49203 15589
rect 49694 15580 49700 15592
rect 49752 15580 49758 15632
rect 51626 15620 51632 15632
rect 51184 15592 51632 15620
rect 7653 15555 7711 15561
rect 7653 15521 7665 15555
rect 7699 15552 7711 15555
rect 8570 15552 8576 15564
rect 7699 15524 8576 15552
rect 7699 15521 7711 15524
rect 7653 15515 7711 15521
rect 8570 15512 8576 15524
rect 8628 15512 8634 15564
rect 10410 15512 10416 15564
rect 10468 15552 10474 15564
rect 10873 15555 10931 15561
rect 10873 15552 10885 15555
rect 10468 15524 10885 15552
rect 10468 15512 10474 15524
rect 10873 15521 10885 15524
rect 10919 15521 10931 15555
rect 12158 15552 12164 15564
rect 12119 15524 12164 15552
rect 10873 15515 10931 15521
rect 12158 15512 12164 15524
rect 12216 15512 12222 15564
rect 12345 15555 12403 15561
rect 12345 15521 12357 15555
rect 12391 15521 12403 15555
rect 12345 15515 12403 15521
rect 13633 15555 13691 15561
rect 13633 15521 13645 15555
rect 13679 15521 13691 15555
rect 13814 15552 13820 15564
rect 13775 15524 13820 15552
rect 13633 15515 13691 15521
rect 5500 15456 7512 15484
rect 5500 15444 5506 15456
rect 10318 15444 10324 15496
rect 10376 15484 10382 15496
rect 12360 15484 12388 15515
rect 10376 15456 12388 15484
rect 13648 15484 13676 15515
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 15470 15552 15476 15564
rect 15431 15524 15476 15552
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 16666 15512 16672 15564
rect 16724 15552 16730 15564
rect 16945 15555 17003 15561
rect 16945 15552 16957 15555
rect 16724 15524 16957 15552
rect 16724 15512 16730 15524
rect 16945 15521 16957 15524
rect 16991 15521 17003 15555
rect 17218 15552 17224 15564
rect 17179 15524 17224 15552
rect 16945 15515 17003 15521
rect 17218 15512 17224 15524
rect 17276 15512 17282 15564
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15552 19487 15555
rect 19702 15552 19708 15564
rect 19475 15524 19708 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 19702 15512 19708 15524
rect 19760 15512 19766 15564
rect 22830 15552 22836 15564
rect 22791 15524 22836 15552
rect 22830 15512 22836 15524
rect 22888 15512 22894 15564
rect 23106 15512 23112 15564
rect 23164 15552 23170 15564
rect 23201 15555 23259 15561
rect 23201 15552 23213 15555
rect 23164 15524 23213 15552
rect 23164 15512 23170 15524
rect 23201 15521 23213 15524
rect 23247 15521 23259 15555
rect 23201 15515 23259 15521
rect 24397 15555 24455 15561
rect 24397 15521 24409 15555
rect 24443 15521 24455 15555
rect 24397 15515 24455 15521
rect 13648 15456 15332 15484
rect 10376 15444 10382 15456
rect 15304 15428 15332 15456
rect 22370 15444 22376 15496
rect 22428 15484 22434 15496
rect 22741 15487 22799 15493
rect 22741 15484 22753 15487
rect 22428 15456 22753 15484
rect 22428 15444 22434 15456
rect 22741 15453 22753 15456
rect 22787 15453 22799 15487
rect 23290 15484 23296 15496
rect 23251 15456 23296 15484
rect 22741 15447 22799 15453
rect 23290 15444 23296 15456
rect 23348 15444 23354 15496
rect 24412 15484 24440 15515
rect 24486 15512 24492 15564
rect 24544 15552 24550 15564
rect 27062 15552 27068 15564
rect 24544 15524 24589 15552
rect 27023 15524 27068 15552
rect 24544 15512 24550 15524
rect 27062 15512 27068 15524
rect 27120 15512 27126 15564
rect 27522 15512 27528 15564
rect 27580 15552 27586 15564
rect 28626 15552 28632 15564
rect 27580 15524 28632 15552
rect 27580 15512 27586 15524
rect 28626 15512 28632 15524
rect 28684 15512 28690 15564
rect 28810 15512 28816 15564
rect 28868 15552 28874 15564
rect 30929 15555 30987 15561
rect 28868 15524 28913 15552
rect 28868 15512 28874 15524
rect 30929 15521 30941 15555
rect 30975 15552 30987 15555
rect 36170 15552 36176 15564
rect 30975 15524 36176 15552
rect 30975 15521 30987 15524
rect 30929 15515 30987 15521
rect 36170 15512 36176 15524
rect 36228 15512 36234 15564
rect 36357 15555 36415 15561
rect 36357 15521 36369 15555
rect 36403 15552 36415 15555
rect 37734 15552 37740 15564
rect 36403 15524 37740 15552
rect 36403 15521 36415 15524
rect 36357 15515 36415 15521
rect 37734 15512 37740 15524
rect 37792 15512 37798 15564
rect 38378 15552 38384 15564
rect 38339 15524 38384 15552
rect 38378 15512 38384 15524
rect 38436 15512 38442 15564
rect 38565 15555 38623 15561
rect 38565 15521 38577 15555
rect 38611 15552 38623 15555
rect 39022 15552 39028 15564
rect 38611 15524 39028 15552
rect 38611 15521 38623 15524
rect 38565 15515 38623 15521
rect 39022 15512 39028 15524
rect 39080 15512 39086 15564
rect 43717 15555 43775 15561
rect 43717 15521 43729 15555
rect 43763 15552 43775 15555
rect 44174 15552 44180 15564
rect 43763 15524 44180 15552
rect 43763 15521 43775 15524
rect 43717 15515 43775 15521
rect 44174 15512 44180 15524
rect 44232 15512 44238 15564
rect 45278 15552 45284 15564
rect 45239 15524 45284 15552
rect 45278 15512 45284 15524
rect 45336 15512 45342 15564
rect 46934 15512 46940 15564
rect 46992 15552 46998 15564
rect 47581 15555 47639 15561
rect 47581 15552 47593 15555
rect 46992 15524 47593 15552
rect 46992 15512 46998 15524
rect 47581 15521 47593 15524
rect 47627 15521 47639 15555
rect 47581 15515 47639 15521
rect 49234 15512 49240 15564
rect 49292 15552 49298 15564
rect 49292 15524 49337 15552
rect 49292 15512 49298 15524
rect 49602 15512 49608 15564
rect 49660 15552 49666 15564
rect 51184 15561 51212 15592
rect 51626 15580 51632 15592
rect 51684 15620 51690 15632
rect 52638 15620 52644 15632
rect 51684 15592 52644 15620
rect 51684 15580 51690 15592
rect 52638 15580 52644 15592
rect 52696 15580 52702 15632
rect 58710 15620 58716 15632
rect 56060 15592 58716 15620
rect 50985 15555 51043 15561
rect 50985 15552 50997 15555
rect 49660 15524 50997 15552
rect 49660 15512 49666 15524
rect 50985 15521 50997 15524
rect 51031 15521 51043 15555
rect 50985 15515 51043 15521
rect 51169 15555 51227 15561
rect 51169 15521 51181 15555
rect 51215 15521 51227 15555
rect 52365 15555 52423 15561
rect 52365 15552 52377 15555
rect 51169 15515 51227 15521
rect 51368 15524 52377 15552
rect 25498 15484 25504 15496
rect 24412 15456 25504 15484
rect 25498 15444 25504 15456
rect 25556 15444 25562 15496
rect 32858 15484 32864 15496
rect 32819 15456 32864 15484
rect 32858 15444 32864 15456
rect 32916 15444 32922 15496
rect 33134 15484 33140 15496
rect 33095 15456 33140 15484
rect 33134 15444 33140 15456
rect 33192 15444 33198 15496
rect 36078 15484 36084 15496
rect 36039 15456 36084 15484
rect 36078 15444 36084 15456
rect 36136 15444 36142 15496
rect 51000 15484 51028 15515
rect 51368 15484 51396 15524
rect 52365 15521 52377 15524
rect 52411 15521 52423 15555
rect 52365 15515 52423 15521
rect 52549 15555 52607 15561
rect 52549 15521 52561 15555
rect 52595 15552 52607 15555
rect 53282 15552 53288 15564
rect 52595 15524 53288 15552
rect 52595 15521 52607 15524
rect 52549 15515 52607 15521
rect 51534 15484 51540 15496
rect 51000 15456 51396 15484
rect 51495 15456 51540 15484
rect 51534 15444 51540 15456
rect 51592 15444 51598 15496
rect 15286 15376 15292 15428
rect 15344 15416 15350 15428
rect 15657 15419 15715 15425
rect 15657 15416 15669 15419
rect 15344 15388 15669 15416
rect 15344 15376 15350 15388
rect 15657 15385 15669 15388
rect 15703 15385 15715 15419
rect 15657 15379 15715 15385
rect 23658 15376 23664 15428
rect 23716 15416 23722 15428
rect 24213 15419 24271 15425
rect 24213 15416 24225 15419
rect 23716 15388 24225 15416
rect 23716 15376 23722 15388
rect 24213 15385 24225 15388
rect 24259 15385 24271 15419
rect 27246 15416 27252 15428
rect 27207 15388 27252 15416
rect 24213 15379 24271 15385
rect 27246 15376 27252 15388
rect 27304 15376 27310 15428
rect 27890 15376 27896 15428
rect 27948 15416 27954 15428
rect 28537 15419 28595 15425
rect 28537 15416 28549 15419
rect 27948 15388 28549 15416
rect 27948 15376 27954 15388
rect 28537 15385 28549 15388
rect 28583 15385 28595 15419
rect 28537 15379 28595 15385
rect 33870 15376 33876 15428
rect 33928 15416 33934 15428
rect 42058 15416 42064 15428
rect 33928 15388 42064 15416
rect 33928 15376 33934 15388
rect 42058 15376 42064 15388
rect 42116 15376 42122 15428
rect 43441 15419 43499 15425
rect 43441 15385 43453 15419
rect 43487 15416 43499 15419
rect 43530 15416 43536 15428
rect 43487 15388 43536 15416
rect 43487 15385 43499 15388
rect 43441 15379 43499 15385
rect 43530 15376 43536 15388
rect 43588 15416 43594 15428
rect 52380 15416 52408 15515
rect 53282 15512 53288 15524
rect 53340 15512 53346 15564
rect 56060 15561 56088 15592
rect 58710 15580 58716 15592
rect 58768 15620 58774 15632
rect 60366 15620 60372 15632
rect 58768 15592 60372 15620
rect 58768 15580 58774 15592
rect 60366 15580 60372 15592
rect 60424 15580 60430 15632
rect 55861 15555 55919 15561
rect 55861 15521 55873 15555
rect 55907 15521 55919 15555
rect 55861 15515 55919 15521
rect 56045 15555 56103 15561
rect 56045 15521 56057 15555
rect 56091 15521 56103 15555
rect 56045 15515 56103 15521
rect 52914 15484 52920 15496
rect 52875 15456 52920 15484
rect 52914 15444 52920 15456
rect 52972 15444 52978 15496
rect 54662 15416 54668 15428
rect 43588 15388 44128 15416
rect 52380 15388 54668 15416
rect 43588 15376 43594 15388
rect 44100 15360 44128 15388
rect 54662 15376 54668 15388
rect 54720 15416 54726 15428
rect 55122 15416 55128 15428
rect 54720 15388 55128 15416
rect 54720 15376 54726 15388
rect 55122 15376 55128 15388
rect 55180 15416 55186 15428
rect 55876 15416 55904 15515
rect 55180 15388 55904 15416
rect 55180 15376 55186 15388
rect 5350 15308 5356 15360
rect 5408 15348 5414 15360
rect 5813 15351 5871 15357
rect 5813 15348 5825 15351
rect 5408 15320 5825 15348
rect 5408 15308 5414 15320
rect 5813 15317 5825 15320
rect 5859 15317 5871 15351
rect 5813 15311 5871 15317
rect 7006 15308 7012 15360
rect 7064 15348 7070 15360
rect 7745 15351 7803 15357
rect 7745 15348 7757 15351
rect 7064 15320 7757 15348
rect 7064 15308 7070 15320
rect 7745 15317 7757 15320
rect 7791 15317 7803 15351
rect 11054 15348 11060 15360
rect 11015 15320 11060 15348
rect 7745 15311 7803 15317
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 12526 15348 12532 15360
rect 12487 15320 12532 15348
rect 12526 15308 12532 15320
rect 12584 15308 12590 15360
rect 19610 15348 19616 15360
rect 19571 15320 19616 15348
rect 19610 15308 19616 15320
rect 19668 15308 19674 15360
rect 22097 15351 22155 15357
rect 22097 15317 22109 15351
rect 22143 15348 22155 15351
rect 27522 15348 27528 15360
rect 22143 15320 27528 15348
rect 22143 15317 22155 15320
rect 22097 15311 22155 15317
rect 27522 15308 27528 15320
rect 27580 15308 27586 15360
rect 31110 15348 31116 15360
rect 31071 15320 31116 15348
rect 31110 15308 31116 15320
rect 31168 15308 31174 15360
rect 33042 15308 33048 15360
rect 33100 15348 33106 15360
rect 34241 15351 34299 15357
rect 34241 15348 34253 15351
rect 33100 15320 34253 15348
rect 33100 15308 33106 15320
rect 34241 15317 34253 15320
rect 34287 15317 34299 15351
rect 36538 15348 36544 15360
rect 36499 15320 36544 15348
rect 34241 15311 34299 15317
rect 36538 15308 36544 15320
rect 36596 15308 36602 15360
rect 38746 15348 38752 15360
rect 38707 15320 38752 15348
rect 38746 15308 38752 15320
rect 38804 15308 38810 15360
rect 43714 15308 43720 15360
rect 43772 15348 43778 15360
rect 43901 15351 43959 15357
rect 43901 15348 43913 15351
rect 43772 15320 43913 15348
rect 43772 15308 43778 15320
rect 43901 15317 43913 15320
rect 43947 15317 43959 15351
rect 43901 15311 43959 15317
rect 44082 15308 44088 15360
rect 44140 15348 44146 15360
rect 45005 15351 45063 15357
rect 45005 15348 45017 15351
rect 44140 15320 45017 15348
rect 44140 15308 44146 15320
rect 45005 15317 45017 15320
rect 45051 15348 45063 15351
rect 47305 15351 47363 15357
rect 47305 15348 47317 15351
rect 45051 15320 47317 15348
rect 45051 15317 45063 15320
rect 45005 15311 45063 15317
rect 47305 15317 47317 15320
rect 47351 15348 47363 15351
rect 48961 15351 49019 15357
rect 48961 15348 48973 15351
rect 47351 15320 48973 15348
rect 47351 15317 47363 15320
rect 47305 15311 47363 15317
rect 48961 15317 48973 15320
rect 49007 15317 49019 15351
rect 48961 15311 49019 15317
rect 53282 15308 53288 15360
rect 53340 15348 53346 15360
rect 54570 15348 54576 15360
rect 53340 15320 54576 15348
rect 53340 15308 53346 15320
rect 54570 15308 54576 15320
rect 54628 15308 54634 15360
rect 55490 15308 55496 15360
rect 55548 15348 55554 15360
rect 56137 15351 56195 15357
rect 56137 15348 56149 15351
rect 55548 15320 56149 15348
rect 55548 15308 55554 15320
rect 56137 15317 56149 15320
rect 56183 15317 56195 15351
rect 56137 15311 56195 15317
rect 1104 15258 62192 15280
rect 1104 15206 11163 15258
rect 11215 15206 11227 15258
rect 11279 15206 11291 15258
rect 11343 15206 11355 15258
rect 11407 15206 31526 15258
rect 31578 15206 31590 15258
rect 31642 15206 31654 15258
rect 31706 15206 31718 15258
rect 31770 15206 51888 15258
rect 51940 15206 51952 15258
rect 52004 15206 52016 15258
rect 52068 15206 52080 15258
rect 52132 15206 62192 15258
rect 1104 15184 62192 15206
rect 8570 15144 8576 15156
rect 8531 15116 8576 15144
rect 8570 15104 8576 15116
rect 8628 15104 8634 15156
rect 15381 15147 15439 15153
rect 15381 15113 15393 15147
rect 15427 15144 15439 15147
rect 16298 15144 16304 15156
rect 15427 15116 16304 15144
rect 15427 15113 15439 15116
rect 15381 15107 15439 15113
rect 16298 15104 16304 15116
rect 16356 15104 16362 15156
rect 16761 15147 16819 15153
rect 16761 15113 16773 15147
rect 16807 15144 16819 15147
rect 16942 15144 16948 15156
rect 16807 15116 16948 15144
rect 16807 15113 16819 15116
rect 16761 15107 16819 15113
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 23014 15104 23020 15156
rect 23072 15144 23078 15156
rect 24121 15147 24179 15153
rect 24121 15144 24133 15147
rect 23072 15116 24133 15144
rect 23072 15104 23078 15116
rect 24121 15113 24133 15116
rect 24167 15113 24179 15147
rect 25498 15144 25504 15156
rect 25459 15116 25504 15144
rect 24121 15107 24179 15113
rect 25498 15104 25504 15116
rect 25556 15104 25562 15156
rect 27890 15104 27896 15156
rect 27948 15144 27954 15156
rect 27985 15147 28043 15153
rect 27985 15144 27997 15147
rect 27948 15116 27997 15144
rect 27948 15104 27954 15116
rect 27985 15113 27997 15116
rect 28031 15113 28043 15147
rect 27985 15107 28043 15113
rect 28626 15104 28632 15156
rect 28684 15144 28690 15156
rect 33042 15144 33048 15156
rect 28684 15116 33048 15144
rect 28684 15104 28690 15116
rect 33042 15104 33048 15116
rect 33100 15104 33106 15156
rect 33134 15104 33140 15156
rect 33192 15144 33198 15156
rect 33689 15147 33747 15153
rect 33689 15144 33701 15147
rect 33192 15116 33701 15144
rect 33192 15104 33198 15116
rect 33689 15113 33701 15116
rect 33735 15113 33747 15147
rect 33689 15107 33747 15113
rect 35158 15104 35164 15156
rect 35216 15144 35222 15156
rect 35621 15147 35679 15153
rect 35621 15144 35633 15147
rect 35216 15116 35633 15144
rect 35216 15104 35222 15116
rect 35621 15113 35633 15116
rect 35667 15113 35679 15147
rect 35621 15107 35679 15113
rect 37366 15104 37372 15156
rect 37424 15144 37430 15156
rect 39025 15147 39083 15153
rect 39025 15144 39037 15147
rect 37424 15116 39037 15144
rect 37424 15104 37430 15116
rect 39025 15113 39037 15116
rect 39071 15113 39083 15147
rect 43530 15144 43536 15156
rect 43491 15116 43536 15144
rect 39025 15107 39083 15113
rect 43530 15104 43536 15116
rect 43588 15104 43594 15156
rect 44450 15104 44456 15156
rect 44508 15144 44514 15156
rect 44729 15147 44787 15153
rect 44729 15144 44741 15147
rect 44508 15116 44741 15144
rect 44508 15104 44514 15116
rect 44729 15113 44741 15116
rect 44775 15113 44787 15147
rect 44729 15107 44787 15113
rect 47673 15147 47731 15153
rect 47673 15113 47685 15147
rect 47719 15144 47731 15147
rect 49602 15144 49608 15156
rect 47719 15116 49608 15144
rect 47719 15113 47731 15116
rect 47673 15107 47731 15113
rect 49602 15104 49608 15116
rect 49660 15104 49666 15156
rect 53282 15144 53288 15156
rect 53243 15116 53288 15144
rect 53282 15104 53288 15116
rect 53340 15104 53346 15156
rect 55401 15147 55459 15153
rect 55401 15113 55413 15147
rect 55447 15144 55459 15147
rect 55582 15144 55588 15156
rect 55447 15116 55588 15144
rect 55447 15113 55459 15116
rect 55401 15107 55459 15113
rect 55582 15104 55588 15116
rect 55640 15104 55646 15156
rect 12434 15036 12440 15088
rect 12492 15036 12498 15088
rect 22480 15048 27844 15076
rect 12452 15008 12480 15036
rect 13817 15011 13875 15017
rect 13817 15008 13829 15011
rect 11164 14980 13829 15008
rect 5353 14943 5411 14949
rect 5353 14909 5365 14943
rect 5399 14940 5411 14943
rect 5442 14940 5448 14952
rect 5399 14912 5448 14940
rect 5399 14909 5411 14912
rect 5353 14903 5411 14909
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 5537 14943 5595 14949
rect 5537 14909 5549 14943
rect 5583 14940 5595 14943
rect 6638 14940 6644 14952
rect 5583 14912 6644 14940
rect 5583 14909 5595 14912
rect 5537 14903 5595 14909
rect 6638 14900 6644 14912
rect 6696 14900 6702 14952
rect 7009 14943 7067 14949
rect 7009 14909 7021 14943
rect 7055 14940 7067 14943
rect 7098 14940 7104 14952
rect 7055 14912 7104 14940
rect 7055 14909 7067 14912
rect 7009 14903 7067 14909
rect 7098 14900 7104 14912
rect 7156 14900 7162 14952
rect 7285 14943 7343 14949
rect 7285 14909 7297 14943
rect 7331 14940 7343 14943
rect 7558 14940 7564 14952
rect 7331 14912 7564 14940
rect 7331 14909 7343 14912
rect 7285 14903 7343 14909
rect 7558 14900 7564 14912
rect 7616 14900 7622 14952
rect 11164 14949 11192 14980
rect 13817 14977 13829 14980
rect 13863 14977 13875 15011
rect 22480 15008 22508 15048
rect 22738 15008 22744 15020
rect 13817 14971 13875 14977
rect 15212 14980 22508 15008
rect 22572 14980 22744 15008
rect 11149 14943 11207 14949
rect 11149 14909 11161 14943
rect 11195 14909 11207 14943
rect 11149 14903 11207 14909
rect 11698 14900 11704 14952
rect 11756 14940 11762 14952
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 11756 14912 12449 14940
rect 11756 14900 11762 14912
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12710 14940 12716 14952
rect 12671 14912 12716 14940
rect 12437 14903 12495 14909
rect 12710 14900 12716 14912
rect 12768 14900 12774 14952
rect 15212 14949 15240 14980
rect 15197 14943 15255 14949
rect 15197 14940 15209 14943
rect 13372 14912 15209 14940
rect 10962 14872 10968 14884
rect 10923 14844 10968 14872
rect 10962 14832 10968 14844
rect 11020 14832 11026 14884
rect 11517 14875 11575 14881
rect 11517 14841 11529 14875
rect 11563 14872 11575 14875
rect 12526 14872 12532 14884
rect 11563 14844 12532 14872
rect 11563 14841 11575 14844
rect 11517 14835 11575 14841
rect 12526 14832 12532 14844
rect 12584 14832 12590 14884
rect 5626 14804 5632 14816
rect 5587 14776 5632 14804
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 10410 14764 10416 14816
rect 10468 14804 10474 14816
rect 13372 14804 13400 14912
rect 15197 14909 15209 14912
rect 15243 14909 15255 14943
rect 16482 14940 16488 14952
rect 16443 14912 16488 14940
rect 15197 14903 15255 14909
rect 16482 14900 16488 14912
rect 16540 14900 16546 14952
rect 16574 14900 16580 14952
rect 16632 14940 16638 14952
rect 16632 14912 16677 14940
rect 16632 14900 16638 14912
rect 18414 14900 18420 14952
rect 18472 14940 18478 14952
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18472 14912 18521 14940
rect 18472 14900 18478 14912
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 18782 14940 18788 14952
rect 18743 14912 18788 14940
rect 18509 14903 18567 14909
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 21174 14900 21180 14952
rect 21232 14940 21238 14952
rect 22189 14943 22247 14949
rect 22189 14940 22201 14943
rect 21232 14912 22201 14940
rect 21232 14900 21238 14912
rect 22189 14909 22201 14912
rect 22235 14909 22247 14943
rect 22189 14903 22247 14909
rect 22281 14943 22339 14949
rect 22281 14909 22293 14943
rect 22327 14940 22339 14943
rect 22370 14940 22376 14952
rect 22327 14912 22376 14940
rect 22327 14909 22339 14912
rect 22281 14903 22339 14909
rect 22370 14900 22376 14912
rect 22428 14900 22434 14952
rect 22572 14949 22600 14980
rect 22738 14968 22744 14980
rect 22796 14968 22802 15020
rect 23658 15008 23664 15020
rect 23619 14980 23664 15008
rect 23658 14968 23664 14980
rect 23716 14968 23722 15020
rect 27816 15008 27844 15048
rect 28166 15036 28172 15088
rect 28224 15076 28230 15088
rect 28224 15048 33548 15076
rect 28224 15036 28230 15048
rect 27816 14980 32168 15008
rect 22557 14943 22615 14949
rect 22557 14909 22569 14943
rect 22603 14909 22615 14943
rect 22557 14903 22615 14909
rect 22649 14943 22707 14949
rect 22649 14909 22661 14943
rect 22695 14940 22707 14943
rect 23014 14940 23020 14952
rect 22695 14912 23020 14940
rect 22695 14909 22707 14912
rect 22649 14903 22707 14909
rect 23014 14900 23020 14912
rect 23072 14940 23078 14952
rect 23290 14940 23296 14952
rect 23072 14912 23296 14940
rect 23072 14900 23078 14912
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 23937 14943 23995 14949
rect 23937 14940 23949 14943
rect 23768 14912 23949 14940
rect 21545 14875 21603 14881
rect 21545 14841 21557 14875
rect 21591 14872 21603 14875
rect 23768 14872 23796 14912
rect 23937 14909 23949 14912
rect 23983 14909 23995 14943
rect 25406 14940 25412 14952
rect 25367 14912 25412 14940
rect 23937 14903 23995 14909
rect 25406 14900 25412 14912
rect 25464 14900 25470 14952
rect 25498 14900 25504 14952
rect 25556 14940 25562 14952
rect 27816 14949 27844 14980
rect 26789 14943 26847 14949
rect 26789 14940 26801 14943
rect 25556 14912 26801 14940
rect 25556 14900 25562 14912
rect 26789 14909 26801 14912
rect 26835 14909 26847 14943
rect 26789 14903 26847 14909
rect 27801 14943 27859 14949
rect 27801 14909 27813 14943
rect 27847 14909 27859 14943
rect 27801 14903 27859 14909
rect 27890 14900 27896 14952
rect 27948 14940 27954 14952
rect 30926 14940 30932 14952
rect 27948 14912 30932 14940
rect 27948 14900 27954 14912
rect 30926 14900 30932 14912
rect 30984 14900 30990 14952
rect 32140 14949 32168 14980
rect 32125 14943 32183 14949
rect 32125 14909 32137 14943
rect 32171 14940 32183 14943
rect 32858 14940 32864 14952
rect 32171 14912 32864 14940
rect 32171 14909 32183 14912
rect 32125 14903 32183 14909
rect 32858 14900 32864 14912
rect 32916 14900 32922 14952
rect 33318 14940 33324 14952
rect 33279 14912 33324 14940
rect 33318 14900 33324 14912
rect 33376 14900 33382 14952
rect 33520 14949 33548 15048
rect 36170 15036 36176 15088
rect 36228 15076 36234 15088
rect 36228 15048 38884 15076
rect 36228 15036 36234 15048
rect 35161 15011 35219 15017
rect 35161 14977 35173 15011
rect 35207 15008 35219 15011
rect 36078 15008 36084 15020
rect 35207 14980 36084 15008
rect 35207 14977 35219 14980
rect 35161 14971 35219 14977
rect 33505 14943 33563 14949
rect 33505 14909 33517 14943
rect 33551 14909 33563 14943
rect 33505 14903 33563 14909
rect 21591 14844 23796 14872
rect 23845 14875 23903 14881
rect 21591 14841 21603 14844
rect 21545 14835 21603 14841
rect 23845 14841 23857 14875
rect 23891 14841 23903 14875
rect 23845 14835 23903 14841
rect 25225 14875 25283 14881
rect 25225 14841 25237 14875
rect 25271 14872 25283 14875
rect 27246 14872 27252 14884
rect 25271 14844 27252 14872
rect 25271 14841 25283 14844
rect 25225 14835 25283 14841
rect 10468 14776 13400 14804
rect 10468 14764 10474 14776
rect 19426 14764 19432 14816
rect 19484 14804 19490 14816
rect 19794 14804 19800 14816
rect 19484 14776 19800 14804
rect 19484 14764 19490 14776
rect 19794 14764 19800 14776
rect 19852 14804 19858 14816
rect 19889 14807 19947 14813
rect 19889 14804 19901 14807
rect 19852 14776 19901 14804
rect 19852 14764 19858 14776
rect 19889 14773 19901 14776
rect 19935 14773 19947 14807
rect 19889 14767 19947 14773
rect 22922 14764 22928 14816
rect 22980 14804 22986 14816
rect 23860 14804 23888 14835
rect 27246 14832 27252 14844
rect 27304 14832 27310 14884
rect 30742 14872 30748 14884
rect 30703 14844 30748 14872
rect 30742 14832 30748 14844
rect 30800 14832 30806 14884
rect 33410 14872 33416 14884
rect 33371 14844 33416 14872
rect 33410 14832 33416 14844
rect 33468 14832 33474 14884
rect 35176 14872 35204 14971
rect 36078 14968 36084 14980
rect 36136 14968 36142 15020
rect 37366 15008 37372 15020
rect 37327 14980 37372 15008
rect 37366 14968 37372 14980
rect 37424 14968 37430 15020
rect 38856 15008 38884 15048
rect 47026 15008 47032 15020
rect 38856 14980 47032 15008
rect 35342 14940 35348 14952
rect 35303 14912 35348 14940
rect 35342 14900 35348 14912
rect 35400 14900 35406 14952
rect 35437 14943 35495 14949
rect 35437 14909 35449 14943
rect 35483 14940 35495 14943
rect 36170 14940 36176 14952
rect 35483 14912 36176 14940
rect 35483 14909 35495 14912
rect 35437 14903 35495 14909
rect 36170 14900 36176 14912
rect 36228 14900 36234 14952
rect 36630 14900 36636 14952
rect 36688 14940 36694 14952
rect 37461 14943 37519 14949
rect 37461 14940 37473 14943
rect 36688 14912 37473 14940
rect 36688 14900 36694 14912
rect 37461 14909 37473 14912
rect 37507 14909 37519 14943
rect 37461 14903 37519 14909
rect 37829 14943 37887 14949
rect 37829 14909 37841 14943
rect 37875 14909 37887 14943
rect 37829 14903 37887 14909
rect 38013 14943 38071 14949
rect 38013 14909 38025 14943
rect 38059 14940 38071 14943
rect 38654 14940 38660 14952
rect 38059 14912 38660 14940
rect 38059 14909 38071 14912
rect 38013 14903 38071 14909
rect 34532 14844 35204 14872
rect 36817 14875 36875 14881
rect 22980 14776 23888 14804
rect 22980 14764 22986 14776
rect 24026 14764 24032 14816
rect 24084 14804 24090 14816
rect 26881 14807 26939 14813
rect 26881 14804 26893 14807
rect 24084 14776 26893 14804
rect 24084 14764 24090 14776
rect 26881 14773 26893 14776
rect 26927 14804 26939 14807
rect 28810 14804 28816 14816
rect 26927 14776 28816 14804
rect 26927 14773 26939 14776
rect 26881 14767 26939 14773
rect 28810 14764 28816 14776
rect 28868 14764 28874 14816
rect 30650 14764 30656 14816
rect 30708 14804 30714 14816
rect 31021 14807 31079 14813
rect 31021 14804 31033 14807
rect 30708 14776 31033 14804
rect 30708 14764 30714 14776
rect 31021 14773 31033 14776
rect 31067 14773 31079 14807
rect 31021 14767 31079 14773
rect 32309 14807 32367 14813
rect 32309 14773 32321 14807
rect 32355 14804 32367 14807
rect 34532 14804 34560 14844
rect 36817 14841 36829 14875
rect 36863 14841 36875 14875
rect 36817 14835 36875 14841
rect 32355 14776 34560 14804
rect 32355 14773 32367 14776
rect 32309 14767 32367 14773
rect 34606 14764 34612 14816
rect 34664 14804 34670 14816
rect 36832 14804 36860 14835
rect 34664 14776 36860 14804
rect 37844 14804 37872 14903
rect 38654 14900 38660 14912
rect 38712 14900 38718 14952
rect 38856 14949 38884 14980
rect 47026 14968 47032 14980
rect 47084 14968 47090 15020
rect 50246 14968 50252 15020
rect 50304 15008 50310 15020
rect 51721 15011 51779 15017
rect 51721 15008 51733 15011
rect 50304 14980 51733 15008
rect 50304 14968 50310 14980
rect 51721 14977 51733 14980
rect 51767 15008 51779 15011
rect 55306 15008 55312 15020
rect 51767 14980 55312 15008
rect 51767 14977 51779 14980
rect 51721 14971 51779 14977
rect 55306 14968 55312 14980
rect 55364 14968 55370 15020
rect 38841 14943 38899 14949
rect 38841 14909 38853 14943
rect 38887 14909 38899 14943
rect 38841 14903 38899 14909
rect 41598 14900 41604 14952
rect 41656 14940 41662 14952
rect 43349 14943 43407 14949
rect 43349 14940 43361 14943
rect 41656 14912 43361 14940
rect 41656 14900 41662 14912
rect 43349 14909 43361 14912
rect 43395 14940 43407 14943
rect 44358 14940 44364 14952
rect 43395 14912 44364 14940
rect 43395 14909 43407 14912
rect 43349 14903 43407 14909
rect 44358 14900 44364 14912
rect 44416 14900 44422 14952
rect 44637 14943 44695 14949
rect 44637 14909 44649 14943
rect 44683 14940 44695 14943
rect 45002 14940 45008 14952
rect 44683 14912 45008 14940
rect 44683 14909 44695 14912
rect 44637 14903 44695 14909
rect 45002 14900 45008 14912
rect 45060 14900 45066 14952
rect 46293 14943 46351 14949
rect 46293 14909 46305 14943
rect 46339 14940 46351 14943
rect 46658 14940 46664 14952
rect 46339 14912 46664 14940
rect 46339 14909 46351 14912
rect 46293 14903 46351 14909
rect 46658 14900 46664 14912
rect 46716 14900 46722 14952
rect 47489 14943 47547 14949
rect 47489 14909 47501 14943
rect 47535 14909 47547 14943
rect 47489 14903 47547 14909
rect 51997 14943 52055 14949
rect 51997 14909 52009 14943
rect 52043 14940 52055 14943
rect 53466 14940 53472 14952
rect 52043 14912 53472 14940
rect 52043 14909 52055 14912
rect 51997 14903 52055 14909
rect 40954 14872 40960 14884
rect 39040 14844 40960 14872
rect 39040 14804 39068 14844
rect 40954 14832 40960 14844
rect 41012 14832 41018 14884
rect 44453 14875 44511 14881
rect 44453 14841 44465 14875
rect 44499 14872 44511 14875
rect 44726 14872 44732 14884
rect 44499 14844 44732 14872
rect 44499 14841 44511 14844
rect 44453 14835 44511 14841
rect 44726 14832 44732 14844
rect 44784 14832 44790 14884
rect 46109 14875 46167 14881
rect 46109 14841 46121 14875
rect 46155 14872 46167 14875
rect 47504 14872 47532 14903
rect 53466 14900 53472 14912
rect 53524 14900 53530 14952
rect 55030 14940 55036 14952
rect 54991 14912 55036 14940
rect 55030 14900 55036 14912
rect 55088 14900 55094 14952
rect 55214 14940 55220 14952
rect 55175 14912 55220 14940
rect 55214 14900 55220 14912
rect 55272 14900 55278 14952
rect 46155 14844 47532 14872
rect 55125 14875 55183 14881
rect 46155 14841 46167 14844
rect 46109 14835 46167 14841
rect 55125 14841 55137 14875
rect 55171 14872 55183 14875
rect 55858 14872 55864 14884
rect 55171 14844 55864 14872
rect 55171 14841 55183 14844
rect 55125 14835 55183 14841
rect 37844 14776 39068 14804
rect 34664 14764 34670 14776
rect 39114 14764 39120 14816
rect 39172 14804 39178 14816
rect 43530 14804 43536 14816
rect 39172 14776 43536 14804
rect 39172 14764 39178 14776
rect 43530 14764 43536 14776
rect 43588 14804 43594 14816
rect 46124 14804 46152 14835
rect 55858 14832 55864 14844
rect 55916 14832 55922 14884
rect 43588 14776 46152 14804
rect 43588 14764 43594 14776
rect 46290 14764 46296 14816
rect 46348 14804 46354 14816
rect 46385 14807 46443 14813
rect 46385 14804 46397 14807
rect 46348 14776 46397 14804
rect 46348 14764 46354 14776
rect 46385 14773 46397 14776
rect 46431 14773 46443 14807
rect 46385 14767 46443 14773
rect 1104 14714 62192 14736
rect 1104 14662 21344 14714
rect 21396 14662 21408 14714
rect 21460 14662 21472 14714
rect 21524 14662 21536 14714
rect 21588 14662 41707 14714
rect 41759 14662 41771 14714
rect 41823 14662 41835 14714
rect 41887 14662 41899 14714
rect 41951 14662 62192 14714
rect 1104 14640 62192 14662
rect 5994 14600 6000 14612
rect 5955 14572 6000 14600
rect 5994 14560 6000 14572
rect 6052 14560 6058 14612
rect 6638 14560 6644 14612
rect 6696 14600 6702 14612
rect 8481 14603 8539 14609
rect 8481 14600 8493 14603
rect 6696 14572 8493 14600
rect 6696 14560 6702 14572
rect 8481 14569 8493 14572
rect 8527 14569 8539 14603
rect 10962 14600 10968 14612
rect 8481 14563 8539 14569
rect 10336 14572 10968 14600
rect 8110 14492 8116 14544
rect 8168 14532 8174 14544
rect 10336 14541 10364 14572
rect 10962 14560 10968 14572
rect 11020 14600 11026 14612
rect 15473 14603 15531 14609
rect 15473 14600 15485 14603
rect 11020 14572 15485 14600
rect 11020 14560 11026 14572
rect 15473 14569 15485 14572
rect 15519 14569 15531 14603
rect 24854 14600 24860 14612
rect 15473 14563 15531 14569
rect 21652 14572 24860 14600
rect 10321 14535 10379 14541
rect 10321 14532 10333 14535
rect 8168 14504 10333 14532
rect 8168 14492 8174 14504
rect 10321 14501 10333 14504
rect 10367 14501 10379 14535
rect 10321 14495 10379 14501
rect 17954 14492 17960 14544
rect 18012 14532 18018 14544
rect 18325 14535 18383 14541
rect 18325 14532 18337 14535
rect 18012 14504 18337 14532
rect 18012 14492 18018 14504
rect 18325 14501 18337 14504
rect 18371 14532 18383 14535
rect 20714 14532 20720 14544
rect 18371 14504 20720 14532
rect 18371 14501 18383 14504
rect 18325 14495 18383 14501
rect 20714 14492 20720 14504
rect 20772 14492 20778 14544
rect 21652 14541 21680 14572
rect 24854 14560 24860 14572
rect 24912 14560 24918 14612
rect 39114 14600 39120 14612
rect 24964 14572 29592 14600
rect 21637 14535 21695 14541
rect 21637 14501 21649 14535
rect 21683 14501 21695 14535
rect 23661 14535 23719 14541
rect 21637 14495 21695 14501
rect 22572 14504 22784 14532
rect 4617 14467 4675 14473
rect 4617 14433 4629 14467
rect 4663 14464 4675 14467
rect 7098 14464 7104 14476
rect 4663 14436 7104 14464
rect 4663 14433 4675 14436
rect 4617 14427 4675 14433
rect 7098 14424 7104 14436
rect 7156 14464 7162 14476
rect 10502 14464 10508 14476
rect 7156 14436 9628 14464
rect 10463 14436 10508 14464
rect 7156 14424 7162 14436
rect 4893 14399 4951 14405
rect 4893 14365 4905 14399
rect 4939 14396 4951 14399
rect 5534 14396 5540 14408
rect 4939 14368 5540 14396
rect 4939 14365 4951 14368
rect 4893 14359 4951 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 7374 14396 7380 14408
rect 7335 14368 7380 14396
rect 7374 14356 7380 14368
rect 7432 14356 7438 14408
rect 9600 14396 9628 14436
rect 10502 14424 10508 14436
rect 10560 14464 10566 14476
rect 15289 14467 15347 14473
rect 10560 14436 13124 14464
rect 10560 14424 10566 14436
rect 11698 14396 11704 14408
rect 9600 14368 11704 14396
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 11977 14399 12035 14405
rect 11977 14365 11989 14399
rect 12023 14396 12035 14399
rect 12986 14396 12992 14408
rect 12023 14368 12992 14396
rect 12023 14365 12035 14368
rect 11977 14359 12035 14365
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 13096 14405 13124 14436
rect 15289 14433 15301 14467
rect 15335 14464 15347 14467
rect 15470 14464 15476 14476
rect 15335 14436 15476 14464
rect 15335 14433 15347 14436
rect 15289 14427 15347 14433
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 16666 14464 16672 14476
rect 16627 14436 16672 14464
rect 16666 14424 16672 14436
rect 16724 14424 16730 14476
rect 19426 14464 19432 14476
rect 19387 14436 19432 14464
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 19518 14424 19524 14476
rect 19576 14464 19582 14476
rect 19981 14467 20039 14473
rect 19576 14436 19621 14464
rect 19576 14424 19582 14436
rect 19981 14433 19993 14467
rect 20027 14464 20039 14467
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 20027 14436 22293 14464
rect 20027 14433 20039 14436
rect 19981 14427 20039 14433
rect 22281 14433 22293 14436
rect 22327 14433 22339 14467
rect 22281 14427 22339 14433
rect 13081 14399 13139 14405
rect 13081 14365 13093 14399
rect 13127 14365 13139 14399
rect 13081 14359 13139 14365
rect 16945 14399 17003 14405
rect 16945 14365 16957 14399
rect 16991 14396 17003 14399
rect 17126 14396 17132 14408
rect 16991 14368 17132 14396
rect 16991 14365 17003 14368
rect 16945 14359 17003 14365
rect 17126 14356 17132 14368
rect 17184 14356 17190 14408
rect 22370 14396 22376 14408
rect 22283 14368 22376 14396
rect 22370 14356 22376 14368
rect 22428 14396 22434 14408
rect 22572 14396 22600 14504
rect 22649 14467 22707 14473
rect 22649 14433 22661 14467
rect 22695 14433 22707 14467
rect 22756 14464 22784 14504
rect 23661 14501 23673 14535
rect 23707 14532 23719 14535
rect 24486 14532 24492 14544
rect 23707 14504 24492 14532
rect 23707 14501 23719 14504
rect 23661 14495 23719 14501
rect 24486 14492 24492 14504
rect 24544 14492 24550 14544
rect 24964 14532 24992 14572
rect 24596 14504 24992 14532
rect 28813 14535 28871 14541
rect 22756 14436 24256 14464
rect 22649 14427 22707 14433
rect 22428 14368 22600 14396
rect 22428 14356 22434 14368
rect 20162 14288 20168 14340
rect 20220 14328 20226 14340
rect 22664 14328 22692 14427
rect 22741 14399 22799 14405
rect 22741 14365 22753 14399
rect 22787 14365 22799 14399
rect 24228 14396 24256 14436
rect 24302 14424 24308 14476
rect 24360 14464 24366 14476
rect 24360 14436 24405 14464
rect 24360 14424 24366 14436
rect 24397 14399 24455 14405
rect 24397 14396 24409 14399
rect 24228 14368 24409 14396
rect 22741 14359 22799 14365
rect 24397 14365 24409 14368
rect 24443 14396 24455 14399
rect 24596 14396 24624 14504
rect 28813 14501 28825 14535
rect 28859 14532 28871 14535
rect 28902 14532 28908 14544
rect 28859 14504 28908 14532
rect 28859 14501 28871 14504
rect 28813 14495 28871 14501
rect 28902 14492 28908 14504
rect 28960 14492 28966 14544
rect 29564 14532 29592 14572
rect 32968 14572 39120 14600
rect 31110 14532 31116 14544
rect 29564 14504 31116 14532
rect 24670 14424 24676 14476
rect 24728 14464 24734 14476
rect 24728 14436 24773 14464
rect 24728 14424 24734 14436
rect 26602 14424 26608 14476
rect 26660 14464 26666 14476
rect 26697 14467 26755 14473
rect 26697 14464 26709 14467
rect 26660 14436 26709 14464
rect 26660 14424 26666 14436
rect 26697 14433 26709 14436
rect 26743 14433 26755 14467
rect 26697 14427 26755 14433
rect 26786 14424 26792 14476
rect 26844 14464 26850 14476
rect 26881 14467 26939 14473
rect 26881 14464 26893 14467
rect 26844 14436 26893 14464
rect 26844 14424 26850 14436
rect 26881 14433 26893 14436
rect 26927 14464 26939 14467
rect 27890 14464 27896 14476
rect 26927 14436 27896 14464
rect 26927 14433 26939 14436
rect 26881 14427 26939 14433
rect 27890 14424 27896 14436
rect 27948 14424 27954 14476
rect 29454 14464 29460 14476
rect 29415 14436 29460 14464
rect 29454 14424 29460 14436
rect 29512 14424 29518 14476
rect 29564 14473 29592 14504
rect 31110 14492 31116 14504
rect 31168 14492 31174 14544
rect 32968 14541 32996 14572
rect 39114 14560 39120 14572
rect 39172 14560 39178 14612
rect 41598 14600 41604 14612
rect 39224 14572 41604 14600
rect 32953 14535 33011 14541
rect 32953 14501 32965 14535
rect 32999 14501 33011 14535
rect 32953 14495 33011 14501
rect 33042 14492 33048 14544
rect 33100 14532 33106 14544
rect 33100 14504 33180 14532
rect 33100 14492 33106 14504
rect 29549 14467 29607 14473
rect 29549 14433 29561 14467
rect 29595 14433 29607 14467
rect 29549 14427 29607 14433
rect 29825 14467 29883 14473
rect 29825 14433 29837 14467
rect 29871 14433 29883 14467
rect 30834 14464 30840 14476
rect 30795 14436 30840 14464
rect 29825 14427 29883 14433
rect 24443 14368 24624 14396
rect 24765 14399 24823 14405
rect 24443 14365 24455 14368
rect 24397 14359 24455 14365
rect 24765 14365 24777 14399
rect 24811 14396 24823 14399
rect 24811 14368 27108 14396
rect 24811 14365 24823 14368
rect 24765 14359 24823 14365
rect 20220 14300 22692 14328
rect 22756 14328 22784 14359
rect 23014 14328 23020 14340
rect 22756 14300 23020 14328
rect 20220 14288 20226 14300
rect 23014 14288 23020 14300
rect 23072 14328 23078 14340
rect 24780 14328 24808 14359
rect 23072 14300 24808 14328
rect 23072 14288 23078 14300
rect 3510 14220 3516 14272
rect 3568 14260 3574 14272
rect 7282 14260 7288 14272
rect 3568 14232 7288 14260
rect 3568 14220 3574 14232
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 10597 14263 10655 14269
rect 10597 14229 10609 14263
rect 10643 14260 10655 14263
rect 14182 14260 14188 14272
rect 10643 14232 14188 14260
rect 10643 14229 10655 14232
rect 10597 14223 10655 14229
rect 14182 14220 14188 14232
rect 14240 14220 14246 14272
rect 22370 14220 22376 14272
rect 22428 14260 22434 14272
rect 26973 14263 27031 14269
rect 26973 14260 26985 14263
rect 22428 14232 26985 14260
rect 22428 14220 22434 14232
rect 26973 14229 26985 14232
rect 27019 14229 27031 14263
rect 27080 14260 27108 14368
rect 28902 14288 28908 14340
rect 28960 14328 28966 14340
rect 29840 14328 29868 14427
rect 30834 14424 30840 14436
rect 30892 14464 30898 14476
rect 33152 14473 33180 14504
rect 33410 14492 33416 14544
rect 33468 14532 33474 14544
rect 33505 14535 33563 14541
rect 33505 14532 33517 14535
rect 33468 14504 33517 14532
rect 33468 14492 33474 14504
rect 33505 14501 33517 14504
rect 33551 14501 33563 14535
rect 33505 14495 33563 14501
rect 34238 14492 34244 14544
rect 34296 14532 34302 14544
rect 34517 14535 34575 14541
rect 34517 14532 34529 14535
rect 34296 14504 34529 14532
rect 34296 14492 34302 14504
rect 34517 14501 34529 14504
rect 34563 14501 34575 14535
rect 34517 14495 34575 14501
rect 35897 14535 35955 14541
rect 35897 14501 35909 14535
rect 35943 14532 35955 14535
rect 37182 14532 37188 14544
rect 35943 14504 37188 14532
rect 35943 14501 35955 14504
rect 35897 14495 35955 14501
rect 37182 14492 37188 14504
rect 37240 14492 37246 14544
rect 39022 14532 39028 14544
rect 38983 14504 39028 14532
rect 39022 14492 39028 14504
rect 39080 14492 39086 14544
rect 33137 14467 33195 14473
rect 30892 14436 33088 14464
rect 30892 14424 30898 14436
rect 29917 14399 29975 14405
rect 29917 14365 29929 14399
rect 29963 14396 29975 14399
rect 33060 14396 33088 14436
rect 33137 14433 33149 14467
rect 33183 14433 33195 14467
rect 34606 14464 34612 14476
rect 34567 14436 34612 14464
rect 33137 14427 33195 14433
rect 34606 14424 34612 14436
rect 34664 14424 34670 14476
rect 35710 14424 35716 14476
rect 35768 14464 35774 14476
rect 36081 14467 36139 14473
rect 36081 14464 36093 14467
rect 35768 14436 36093 14464
rect 35768 14424 35774 14436
rect 36081 14433 36093 14436
rect 36127 14433 36139 14467
rect 37909 14467 37967 14473
rect 37909 14464 37921 14467
rect 36081 14427 36139 14433
rect 37660 14436 37921 14464
rect 37660 14408 37688 14436
rect 37909 14433 37921 14436
rect 37955 14433 37967 14467
rect 37909 14427 37967 14433
rect 38562 14424 38568 14476
rect 38620 14464 38626 14476
rect 39224 14464 39252 14572
rect 41598 14560 41604 14572
rect 41656 14560 41662 14612
rect 42058 14560 42064 14612
rect 42116 14600 42122 14612
rect 43809 14603 43867 14609
rect 43809 14600 43821 14603
rect 42116 14572 43821 14600
rect 42116 14560 42122 14572
rect 43809 14569 43821 14572
rect 43855 14569 43867 14603
rect 47210 14600 47216 14612
rect 43809 14563 43867 14569
rect 44836 14572 47216 14600
rect 43714 14492 43720 14544
rect 43772 14532 43778 14544
rect 44836 14532 44864 14572
rect 47210 14560 47216 14572
rect 47268 14560 47274 14612
rect 51626 14600 51632 14612
rect 51587 14572 51632 14600
rect 51626 14560 51632 14572
rect 51684 14560 51690 14612
rect 43772 14504 44864 14532
rect 46385 14535 46443 14541
rect 43772 14492 43778 14504
rect 46385 14501 46397 14535
rect 46431 14532 46443 14535
rect 46658 14532 46664 14544
rect 46431 14504 46664 14532
rect 46431 14501 46443 14504
rect 46385 14495 46443 14501
rect 46658 14492 46664 14504
rect 46716 14492 46722 14544
rect 52914 14532 52920 14544
rect 52875 14504 52920 14532
rect 52914 14492 52920 14504
rect 52972 14492 52978 14544
rect 53466 14532 53472 14544
rect 53427 14504 53472 14532
rect 53466 14492 53472 14504
rect 53524 14492 53530 14544
rect 56229 14535 56287 14541
rect 56229 14501 56241 14535
rect 56275 14532 56287 14535
rect 56502 14532 56508 14544
rect 56275 14504 56508 14532
rect 56275 14501 56287 14504
rect 56229 14495 56287 14501
rect 56502 14492 56508 14504
rect 56560 14492 56566 14544
rect 58710 14532 58716 14544
rect 58671 14504 58716 14532
rect 58710 14492 58716 14504
rect 58768 14492 58774 14544
rect 38620 14436 39252 14464
rect 39669 14467 39727 14473
rect 38620 14424 38626 14436
rect 39669 14433 39681 14467
rect 39715 14433 39727 14467
rect 39669 14427 39727 14433
rect 40037 14467 40095 14473
rect 40037 14433 40049 14467
rect 40083 14464 40095 14467
rect 43622 14464 43628 14476
rect 40083 14436 41460 14464
rect 43583 14436 43628 14464
rect 40083 14433 40095 14436
rect 40037 14427 40095 14433
rect 37642 14396 37648 14408
rect 29963 14368 31064 14396
rect 33060 14368 37648 14396
rect 29963 14365 29975 14368
rect 29917 14359 29975 14365
rect 28960 14300 29868 14328
rect 28960 14288 28966 14300
rect 29932 14260 29960 14359
rect 31036 14337 31064 14368
rect 37642 14356 37648 14368
rect 37700 14356 37706 14408
rect 38470 14356 38476 14408
rect 38528 14396 38534 14408
rect 39577 14399 39635 14405
rect 39577 14396 39589 14399
rect 38528 14368 39589 14396
rect 38528 14356 38534 14368
rect 39577 14365 39589 14368
rect 39623 14365 39635 14399
rect 39577 14359 39635 14365
rect 31021 14331 31079 14337
rect 31021 14297 31033 14331
rect 31067 14297 31079 14331
rect 31021 14291 31079 14297
rect 34333 14331 34391 14337
rect 34333 14297 34345 14331
rect 34379 14328 34391 14331
rect 36078 14328 36084 14340
rect 34379 14300 36084 14328
rect 34379 14297 34391 14300
rect 34333 14291 34391 14297
rect 36078 14288 36084 14300
rect 36136 14288 36142 14340
rect 38105 14331 38163 14337
rect 38105 14297 38117 14331
rect 38151 14328 38163 14331
rect 38654 14328 38660 14340
rect 38151 14300 38660 14328
rect 38151 14297 38163 14300
rect 38105 14291 38163 14297
rect 38654 14288 38660 14300
rect 38712 14328 38718 14340
rect 39390 14328 39396 14340
rect 38712 14300 39396 14328
rect 38712 14288 38718 14300
rect 39390 14288 39396 14300
rect 39448 14288 39454 14340
rect 39684 14328 39712 14427
rect 39850 14356 39856 14408
rect 39908 14396 39914 14408
rect 40129 14399 40187 14405
rect 40129 14396 40141 14399
rect 39908 14368 40141 14396
rect 39908 14356 39914 14368
rect 40129 14365 40141 14368
rect 40175 14365 40187 14399
rect 41432 14396 41460 14436
rect 43622 14424 43628 14436
rect 43680 14424 43686 14476
rect 44729 14467 44787 14473
rect 44729 14433 44741 14467
rect 44775 14464 44787 14467
rect 45922 14464 45928 14476
rect 44775 14436 45928 14464
rect 44775 14433 44787 14436
rect 44729 14427 44787 14433
rect 45922 14424 45928 14436
rect 45980 14424 45986 14476
rect 46106 14424 46112 14476
rect 46164 14464 46170 14476
rect 47213 14467 47271 14473
rect 47213 14464 47225 14467
rect 46164 14436 47225 14464
rect 46164 14424 46170 14436
rect 47213 14433 47225 14436
rect 47259 14433 47271 14467
rect 47213 14427 47271 14433
rect 48038 14424 48044 14476
rect 48096 14464 48102 14476
rect 50246 14464 50252 14476
rect 48096 14436 50252 14464
rect 48096 14424 48102 14436
rect 50246 14424 50252 14436
rect 50304 14424 50310 14476
rect 53006 14464 53012 14476
rect 52967 14436 53012 14464
rect 53006 14424 53012 14436
rect 53064 14424 53070 14476
rect 54573 14467 54631 14473
rect 54573 14433 54585 14467
rect 54619 14464 54631 14467
rect 55306 14464 55312 14476
rect 54619 14436 55312 14464
rect 54619 14433 54631 14436
rect 54573 14427 54631 14433
rect 55306 14424 55312 14436
rect 55364 14464 55370 14476
rect 55364 14436 56456 14464
rect 55364 14424 55370 14436
rect 56428 14408 56456 14436
rect 44450 14396 44456 14408
rect 41432 14368 44456 14396
rect 40129 14359 40187 14365
rect 44450 14356 44456 14368
rect 44508 14356 44514 14408
rect 45005 14399 45063 14405
rect 45005 14365 45017 14399
rect 45051 14396 45063 14399
rect 46566 14396 46572 14408
rect 45051 14368 46572 14396
rect 45051 14365 45063 14368
rect 45005 14359 45063 14365
rect 46566 14356 46572 14368
rect 46624 14356 46630 14408
rect 50525 14399 50583 14405
rect 50525 14365 50537 14399
rect 50571 14396 50583 14399
rect 52178 14396 52184 14408
rect 50571 14368 52184 14396
rect 50571 14365 50583 14368
rect 50525 14359 50583 14365
rect 52178 14356 52184 14368
rect 52236 14356 52242 14408
rect 54846 14396 54852 14408
rect 54807 14368 54852 14396
rect 54846 14356 54852 14368
rect 54904 14356 54910 14408
rect 56410 14356 56416 14408
rect 56468 14396 56474 14408
rect 57057 14399 57115 14405
rect 57057 14396 57069 14399
rect 56468 14368 57069 14396
rect 56468 14356 56474 14368
rect 57057 14365 57069 14368
rect 57103 14365 57115 14399
rect 57330 14396 57336 14408
rect 57291 14368 57336 14396
rect 57057 14359 57115 14365
rect 57330 14356 57336 14368
rect 57388 14356 57394 14408
rect 40770 14328 40776 14340
rect 39684 14300 40776 14328
rect 40770 14288 40776 14300
rect 40828 14288 40834 14340
rect 27080 14232 29960 14260
rect 26973 14223 27031 14229
rect 30926 14220 30932 14272
rect 30984 14260 30990 14272
rect 32490 14260 32496 14272
rect 30984 14232 32496 14260
rect 30984 14220 30990 14232
rect 32490 14220 32496 14232
rect 32548 14220 32554 14272
rect 34790 14260 34796 14272
rect 34751 14232 34796 14260
rect 34790 14220 34796 14232
rect 34848 14220 34854 14272
rect 34882 14220 34888 14272
rect 34940 14260 34946 14272
rect 36173 14263 36231 14269
rect 36173 14260 36185 14263
rect 34940 14232 36185 14260
rect 34940 14220 34946 14232
rect 36173 14229 36185 14232
rect 36219 14229 36231 14263
rect 36173 14223 36231 14229
rect 39114 14220 39120 14272
rect 39172 14260 39178 14272
rect 45462 14260 45468 14272
rect 39172 14232 45468 14260
rect 39172 14220 39178 14232
rect 45462 14220 45468 14232
rect 45520 14220 45526 14272
rect 47397 14263 47455 14269
rect 47397 14229 47409 14263
rect 47443 14260 47455 14263
rect 52730 14260 52736 14272
rect 47443 14232 52736 14260
rect 47443 14229 47455 14232
rect 47397 14223 47455 14229
rect 52730 14220 52736 14232
rect 52788 14220 52794 14272
rect 1104 14170 62192 14192
rect 1104 14118 11163 14170
rect 11215 14118 11227 14170
rect 11279 14118 11291 14170
rect 11343 14118 11355 14170
rect 11407 14118 31526 14170
rect 31578 14118 31590 14170
rect 31642 14118 31654 14170
rect 31706 14118 31718 14170
rect 31770 14118 51888 14170
rect 51940 14118 51952 14170
rect 52004 14118 52016 14170
rect 52068 14118 52080 14170
rect 52132 14118 62192 14170
rect 1104 14096 62192 14118
rect 5258 14016 5264 14068
rect 5316 14056 5322 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 5316 14028 6837 14056
rect 5316 14016 5322 14028
rect 6825 14025 6837 14028
rect 6871 14056 6883 14059
rect 11054 14056 11060 14068
rect 6871 14028 11060 14056
rect 6871 14025 6883 14028
rect 6825 14019 6883 14025
rect 11054 14016 11060 14028
rect 11112 14056 11118 14068
rect 12342 14056 12348 14068
rect 11112 14028 12348 14056
rect 11112 14016 11118 14028
rect 12342 14016 12348 14028
rect 12400 14056 12406 14068
rect 12437 14059 12495 14065
rect 12437 14056 12449 14059
rect 12400 14028 12449 14056
rect 12400 14016 12406 14028
rect 12437 14025 12449 14028
rect 12483 14025 12495 14059
rect 12437 14019 12495 14025
rect 12710 14016 12716 14068
rect 12768 14056 12774 14068
rect 12897 14059 12955 14065
rect 12897 14056 12909 14059
rect 12768 14028 12909 14056
rect 12768 14016 12774 14028
rect 12897 14025 12909 14028
rect 12943 14025 12955 14059
rect 12897 14019 12955 14025
rect 12986 14016 12992 14068
rect 13044 14056 13050 14068
rect 14461 14059 14519 14065
rect 14461 14056 14473 14059
rect 13044 14028 14473 14056
rect 13044 14016 13050 14028
rect 14461 14025 14473 14028
rect 14507 14025 14519 14059
rect 14461 14019 14519 14025
rect 18417 14059 18475 14065
rect 18417 14025 18429 14059
rect 18463 14025 18475 14059
rect 22462 14056 22468 14068
rect 22423 14028 22468 14056
rect 18417 14019 18475 14025
rect 7190 13988 7196 14000
rect 5736 13960 7196 13988
rect 5626 13920 5632 13932
rect 5368 13892 5632 13920
rect 5258 13852 5264 13864
rect 5219 13824 5264 13852
rect 5258 13812 5264 13824
rect 5316 13812 5322 13864
rect 5368 13861 5396 13892
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 5353 13855 5411 13861
rect 5353 13821 5365 13855
rect 5399 13821 5411 13855
rect 5353 13815 5411 13821
rect 5445 13855 5503 13861
rect 5445 13821 5457 13855
rect 5491 13852 5503 13855
rect 5736 13852 5764 13960
rect 7190 13948 7196 13960
rect 7248 13948 7254 14000
rect 7282 13948 7288 14000
rect 7340 13988 7346 14000
rect 18432 13988 18460 14019
rect 22462 14016 22468 14028
rect 22520 14016 22526 14068
rect 24302 14016 24308 14068
rect 24360 14056 24366 14068
rect 24581 14059 24639 14065
rect 24581 14056 24593 14059
rect 24360 14028 24593 14056
rect 24360 14016 24366 14028
rect 24581 14025 24593 14028
rect 24627 14025 24639 14059
rect 29270 14056 29276 14068
rect 24581 14019 24639 14025
rect 25884 14028 29276 14056
rect 7340 13960 18460 13988
rect 7340 13948 7346 13960
rect 24118 13948 24124 14000
rect 24176 13988 24182 14000
rect 25884 13988 25912 14028
rect 29270 14016 29276 14028
rect 29328 14016 29334 14068
rect 29454 14016 29460 14068
rect 29512 14056 29518 14068
rect 32953 14059 33011 14065
rect 32953 14056 32965 14059
rect 29512 14028 32965 14056
rect 29512 14016 29518 14028
rect 32953 14025 32965 14028
rect 32999 14025 33011 14059
rect 32953 14019 33011 14025
rect 33318 14016 33324 14068
rect 33376 14056 33382 14068
rect 35069 14059 35127 14065
rect 35069 14056 35081 14059
rect 33376 14028 35081 14056
rect 33376 14016 33382 14028
rect 35069 14025 35081 14028
rect 35115 14056 35127 14059
rect 38562 14056 38568 14068
rect 35115 14028 38568 14056
rect 35115 14025 35127 14028
rect 35069 14019 35127 14025
rect 38562 14016 38568 14028
rect 38620 14016 38626 14068
rect 44085 14059 44143 14065
rect 44085 14025 44097 14059
rect 44131 14056 44143 14059
rect 44174 14056 44180 14068
rect 44131 14028 44180 14056
rect 44131 14025 44143 14028
rect 44085 14019 44143 14025
rect 44174 14016 44180 14028
rect 44232 14016 44238 14068
rect 44358 14016 44364 14068
rect 44416 14056 44422 14068
rect 46106 14056 46112 14068
rect 44416 14028 46112 14056
rect 44416 14016 44422 14028
rect 46106 14016 46112 14028
rect 46164 14016 46170 14068
rect 46566 14056 46572 14068
rect 46527 14028 46572 14056
rect 46566 14016 46572 14028
rect 46624 14016 46630 14068
rect 52178 14056 52184 14068
rect 52139 14028 52184 14056
rect 52178 14016 52184 14028
rect 52236 14016 52242 14068
rect 52730 14016 52736 14068
rect 52788 14056 52794 14068
rect 53745 14059 53803 14065
rect 53745 14056 53757 14059
rect 52788 14028 53757 14056
rect 52788 14016 52794 14028
rect 53745 14025 53757 14028
rect 53791 14056 53803 14059
rect 55030 14056 55036 14068
rect 53791 14028 55036 14056
rect 53791 14025 53803 14028
rect 53745 14019 53803 14025
rect 55030 14016 55036 14028
rect 55088 14056 55094 14068
rect 55309 14059 55367 14065
rect 55309 14056 55321 14059
rect 55088 14028 55321 14056
rect 55088 14016 55094 14028
rect 55309 14025 55321 14028
rect 55355 14025 55367 14059
rect 55309 14019 55367 14025
rect 37366 13988 37372 14000
rect 24176 13960 25912 13988
rect 24176 13948 24182 13960
rect 25884 13932 25912 13960
rect 36924 13960 37372 13988
rect 5905 13923 5963 13929
rect 5905 13889 5917 13923
rect 5951 13920 5963 13923
rect 7374 13920 7380 13932
rect 5951 13892 7380 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 7558 13920 7564 13932
rect 7519 13892 7564 13920
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 12342 13880 12348 13932
rect 12400 13920 12406 13932
rect 14001 13923 14059 13929
rect 14001 13920 14013 13923
rect 12400 13892 14013 13920
rect 12400 13880 12406 13892
rect 14001 13889 14013 13892
rect 14047 13889 14059 13923
rect 18138 13920 18144 13932
rect 18099 13892 18144 13920
rect 14001 13883 14059 13889
rect 18138 13880 18144 13892
rect 18196 13880 18202 13932
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 19521 13923 19579 13929
rect 19521 13920 19533 13923
rect 18472 13892 19533 13920
rect 18472 13880 18478 13892
rect 19521 13889 19533 13892
rect 19567 13889 19579 13923
rect 19521 13883 19579 13889
rect 23014 13880 23020 13932
rect 23072 13920 23078 13932
rect 25866 13920 25872 13932
rect 23072 13892 24440 13920
rect 25779 13892 25872 13920
rect 23072 13880 23078 13892
rect 5491 13824 5764 13852
rect 5491 13821 5503 13824
rect 5445 13815 5503 13821
rect 5810 13812 5816 13864
rect 5868 13852 5874 13864
rect 7006 13852 7012 13864
rect 5868 13824 6776 13852
rect 6967 13824 7012 13852
rect 5868 13812 5874 13824
rect 6748 13784 6776 13824
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 7101 13855 7159 13861
rect 7101 13821 7113 13855
rect 7147 13821 7159 13855
rect 7101 13815 7159 13821
rect 7116 13784 7144 13815
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 10965 13855 11023 13861
rect 10965 13852 10977 13855
rect 8352 13824 10977 13852
rect 8352 13812 8358 13824
rect 10965 13821 10977 13824
rect 11011 13821 11023 13855
rect 10965 13815 11023 13821
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 11333 13855 11391 13861
rect 11112 13824 11157 13852
rect 11112 13812 11118 13824
rect 11333 13821 11345 13855
rect 11379 13821 11391 13855
rect 11514 13852 11520 13864
rect 11475 13824 11520 13852
rect 11333 13815 11391 13821
rect 10318 13784 10324 13796
rect 6748 13756 7144 13784
rect 10279 13756 10324 13784
rect 10318 13744 10324 13756
rect 10376 13744 10382 13796
rect 11348 13784 11376 13815
rect 11514 13812 11520 13824
rect 11572 13812 11578 13864
rect 12710 13852 12716 13864
rect 12671 13824 12716 13852
rect 12710 13812 12716 13824
rect 12768 13812 12774 13864
rect 13722 13812 13728 13864
rect 13780 13852 13786 13864
rect 14277 13855 14335 13861
rect 14277 13852 14289 13855
rect 13780 13824 14289 13852
rect 13780 13812 13786 13824
rect 14277 13821 14289 13824
rect 14323 13821 14335 13855
rect 18230 13852 18236 13864
rect 18191 13824 18236 13852
rect 14277 13815 14335 13821
rect 18230 13812 18236 13824
rect 18288 13812 18294 13864
rect 19797 13855 19855 13861
rect 19797 13821 19809 13855
rect 19843 13852 19855 13855
rect 20898 13852 20904 13864
rect 19843 13824 20904 13852
rect 19843 13821 19855 13824
rect 19797 13815 19855 13821
rect 20898 13812 20904 13824
rect 20956 13812 20962 13864
rect 22094 13812 22100 13864
rect 22152 13852 22158 13864
rect 22278 13852 22284 13864
rect 22152 13824 22197 13852
rect 22239 13824 22284 13852
rect 22152 13812 22158 13824
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 22370 13812 22376 13864
rect 22428 13812 22434 13864
rect 24412 13861 24440 13892
rect 25866 13880 25872 13892
rect 25924 13880 25930 13932
rect 26602 13920 26608 13932
rect 25976 13892 26608 13920
rect 24305 13855 24363 13861
rect 24305 13821 24317 13855
rect 24351 13821 24363 13855
rect 24305 13815 24363 13821
rect 24397 13855 24455 13861
rect 24397 13821 24409 13855
rect 24443 13821 24455 13855
rect 24397 13815 24455 13821
rect 24596 13824 25820 13852
rect 11698 13784 11704 13796
rect 11348 13756 11704 13784
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 12526 13744 12532 13796
rect 12584 13784 12590 13796
rect 12621 13787 12679 13793
rect 12621 13784 12633 13787
rect 12584 13756 12633 13784
rect 12584 13744 12590 13756
rect 12621 13753 12633 13756
rect 12667 13753 12679 13787
rect 14182 13784 14188 13796
rect 14143 13756 14188 13784
rect 12621 13747 12679 13753
rect 14182 13744 14188 13756
rect 14240 13744 14246 13796
rect 15378 13744 15384 13796
rect 15436 13784 15442 13796
rect 18322 13784 18328 13796
rect 15436 13756 18328 13784
rect 15436 13744 15442 13756
rect 18322 13744 18328 13756
rect 18380 13744 18386 13796
rect 22189 13787 22247 13793
rect 20456 13756 21864 13784
rect 3326 13676 3332 13728
rect 3384 13716 3390 13728
rect 20456 13716 20484 13756
rect 3384 13688 20484 13716
rect 21085 13719 21143 13725
rect 3384 13676 3390 13688
rect 21085 13685 21097 13719
rect 21131 13716 21143 13719
rect 21726 13716 21732 13728
rect 21131 13688 21732 13716
rect 21131 13685 21143 13688
rect 21085 13679 21143 13685
rect 21726 13676 21732 13688
rect 21784 13676 21790 13728
rect 21836 13716 21864 13756
rect 22189 13753 22201 13787
rect 22235 13784 22247 13787
rect 22388 13784 22416 13812
rect 22235 13756 22416 13784
rect 24320 13784 24348 13815
rect 24596 13784 24624 13824
rect 24320 13756 24624 13784
rect 25792 13784 25820 13824
rect 25976 13784 26004 13892
rect 26602 13880 26608 13892
rect 26660 13920 26666 13932
rect 27249 13923 27307 13929
rect 27249 13920 27261 13923
rect 26660 13892 27261 13920
rect 26660 13880 26666 13892
rect 27249 13889 27261 13892
rect 27295 13889 27307 13923
rect 27249 13883 27307 13889
rect 29270 13880 29276 13932
rect 29328 13920 29334 13932
rect 36924 13929 36952 13960
rect 37366 13948 37372 13960
rect 37424 13948 37430 14000
rect 37642 13948 37648 14000
rect 37700 13988 37706 14000
rect 43714 13988 43720 14000
rect 37700 13960 43720 13988
rect 37700 13948 37706 13960
rect 43714 13948 43720 13960
rect 43772 13948 43778 14000
rect 48041 13991 48099 13997
rect 48041 13957 48053 13991
rect 48087 13957 48099 13991
rect 48041 13951 48099 13957
rect 50709 13991 50767 13997
rect 50709 13957 50721 13991
rect 50755 13957 50767 13991
rect 50709 13951 50767 13957
rect 51721 13991 51779 13997
rect 51721 13957 51733 13991
rect 51767 13988 51779 13991
rect 52748 13988 52776 14016
rect 51767 13960 52776 13988
rect 51767 13957 51779 13960
rect 51721 13951 51779 13957
rect 30193 13923 30251 13929
rect 30193 13920 30205 13923
rect 29328 13892 30205 13920
rect 29328 13880 29334 13892
rect 30193 13889 30205 13892
rect 30239 13889 30251 13923
rect 30193 13883 30251 13889
rect 31573 13923 31631 13929
rect 31573 13889 31585 13923
rect 31619 13920 31631 13923
rect 32677 13923 32735 13929
rect 32677 13920 32689 13923
rect 31619 13892 32689 13920
rect 31619 13889 31631 13892
rect 31573 13883 31631 13889
rect 32677 13889 32689 13892
rect 32723 13889 32735 13923
rect 32677 13883 32735 13889
rect 36909 13923 36967 13929
rect 36909 13889 36921 13923
rect 36955 13889 36967 13923
rect 39114 13920 39120 13932
rect 36909 13883 36967 13889
rect 37200 13892 39120 13920
rect 26142 13852 26148 13864
rect 26103 13824 26148 13852
rect 26142 13812 26148 13824
rect 26200 13812 26206 13864
rect 30466 13852 30472 13864
rect 30427 13824 30472 13852
rect 30466 13812 30472 13824
rect 30524 13812 30530 13864
rect 30742 13812 30748 13864
rect 30800 13852 30806 13864
rect 31588 13852 31616 13883
rect 30800 13824 31616 13852
rect 32769 13855 32827 13861
rect 30800 13812 30806 13824
rect 32769 13821 32781 13855
rect 32815 13821 32827 13855
rect 32769 13815 32827 13821
rect 25792 13756 26004 13784
rect 22235 13753 22247 13756
rect 22189 13747 22247 13753
rect 27062 13744 27068 13796
rect 27120 13784 27126 13796
rect 30282 13784 30288 13796
rect 27120 13756 30288 13784
rect 27120 13744 27126 13756
rect 30282 13744 30288 13756
rect 30340 13744 30346 13796
rect 32784 13784 32812 13815
rect 32858 13812 32864 13864
rect 32916 13852 32922 13864
rect 34885 13855 34943 13861
rect 34885 13852 34897 13855
rect 32916 13824 34897 13852
rect 32916 13812 32922 13824
rect 34885 13821 34897 13824
rect 34931 13821 34943 13855
rect 36814 13852 36820 13864
rect 36775 13824 36820 13852
rect 34885 13815 34943 13821
rect 36814 13812 36820 13824
rect 36872 13812 36878 13864
rect 37200 13861 37228 13892
rect 39114 13880 39120 13892
rect 39172 13880 39178 13932
rect 47394 13920 47400 13932
rect 44744 13892 47400 13920
rect 44744 13864 44772 13892
rect 47394 13880 47400 13892
rect 47452 13920 47458 13932
rect 48056 13920 48084 13951
rect 48222 13920 48228 13932
rect 47452 13892 48228 13920
rect 47452 13880 47458 13892
rect 48222 13880 48228 13892
rect 48280 13880 48286 13932
rect 37185 13855 37243 13861
rect 37185 13821 37197 13855
rect 37231 13821 37243 13855
rect 37185 13815 37243 13821
rect 37369 13855 37427 13861
rect 37369 13821 37381 13855
rect 37415 13852 37427 13855
rect 38654 13852 38660 13864
rect 37415 13824 38660 13852
rect 37415 13821 37427 13824
rect 37369 13815 37427 13821
rect 38654 13812 38660 13824
rect 38712 13812 38718 13864
rect 38838 13852 38844 13864
rect 38799 13824 38844 13852
rect 38838 13812 38844 13824
rect 38896 13812 38902 13864
rect 38933 13855 38991 13861
rect 38933 13821 38945 13855
rect 38979 13821 38991 13855
rect 38933 13815 38991 13821
rect 39209 13855 39267 13861
rect 39209 13821 39221 13855
rect 39255 13821 39267 13855
rect 39390 13852 39396 13864
rect 39303 13824 39396 13852
rect 39209 13815 39267 13821
rect 35158 13784 35164 13796
rect 32784 13756 35164 13784
rect 35158 13744 35164 13756
rect 35216 13744 35222 13796
rect 36170 13784 36176 13796
rect 36131 13756 36176 13784
rect 36170 13744 36176 13756
rect 36228 13744 36234 13796
rect 38194 13784 38200 13796
rect 38155 13756 38200 13784
rect 38194 13744 38200 13756
rect 38252 13744 38258 13796
rect 38948 13784 38976 13815
rect 38580 13756 38976 13784
rect 31110 13716 31116 13728
rect 21836 13688 31116 13716
rect 31110 13676 31116 13688
rect 31168 13676 31174 13728
rect 37366 13676 37372 13728
rect 37424 13716 37430 13728
rect 38470 13716 38476 13728
rect 37424 13688 38476 13716
rect 37424 13676 37430 13688
rect 38470 13676 38476 13688
rect 38528 13716 38534 13728
rect 38580 13716 38608 13756
rect 38528 13688 38608 13716
rect 39224 13716 39252 13815
rect 39390 13812 39396 13824
rect 39448 13852 39454 13864
rect 39850 13852 39856 13864
rect 39448 13824 39856 13852
rect 39448 13812 39454 13824
rect 39850 13812 39856 13824
rect 39908 13812 39914 13864
rect 44082 13812 44088 13864
rect 44140 13852 44146 13864
rect 44637 13855 44695 13861
rect 44637 13852 44649 13855
rect 44140 13824 44649 13852
rect 44140 13812 44146 13824
rect 44637 13821 44649 13824
rect 44683 13821 44695 13855
rect 44637 13815 44695 13821
rect 44726 13812 44732 13864
rect 44784 13852 44790 13864
rect 44784 13824 44829 13852
rect 44784 13812 44790 13824
rect 44910 13812 44916 13864
rect 44968 13852 44974 13864
rect 45005 13855 45063 13861
rect 45005 13852 45017 13855
rect 44968 13824 45017 13852
rect 44968 13812 44974 13824
rect 45005 13821 45017 13824
rect 45051 13821 45063 13855
rect 45005 13815 45063 13821
rect 45189 13855 45247 13861
rect 45189 13821 45201 13855
rect 45235 13852 45247 13855
rect 45646 13852 45652 13864
rect 45235 13824 45652 13852
rect 45235 13821 45247 13824
rect 45189 13815 45247 13821
rect 45646 13812 45652 13824
rect 45704 13812 45710 13864
rect 46382 13852 46388 13864
rect 46343 13824 46388 13852
rect 46382 13812 46388 13824
rect 46440 13812 46446 13864
rect 47026 13812 47032 13864
rect 47084 13852 47090 13864
rect 47857 13855 47915 13861
rect 47857 13852 47869 13855
rect 47084 13824 47869 13852
rect 47084 13812 47090 13824
rect 47857 13821 47869 13824
rect 47903 13821 47915 13855
rect 48961 13855 49019 13861
rect 48961 13852 48973 13855
rect 47857 13815 47915 13821
rect 47964 13824 48973 13852
rect 46290 13784 46296 13796
rect 46251 13756 46296 13784
rect 46290 13744 46296 13756
rect 46348 13744 46354 13796
rect 47210 13744 47216 13796
rect 47268 13784 47274 13796
rect 47964 13784 47992 13824
rect 48961 13821 48973 13824
rect 49007 13852 49019 13855
rect 50525 13855 50583 13861
rect 50525 13852 50537 13855
rect 49007 13824 50537 13852
rect 49007 13821 49019 13824
rect 48961 13815 49019 13821
rect 50525 13821 50537 13824
rect 50571 13821 50583 13855
rect 50724 13852 50752 13951
rect 51534 13880 51540 13932
rect 51592 13920 51598 13932
rect 54481 13923 54539 13929
rect 51592 13892 51948 13920
rect 51592 13880 51598 13892
rect 51920 13861 51948 13892
rect 54481 13889 54493 13923
rect 54527 13920 54539 13923
rect 54846 13920 54852 13932
rect 54527 13892 54852 13920
rect 54527 13889 54539 13892
rect 54481 13883 54539 13889
rect 54846 13880 54852 13892
rect 54904 13880 54910 13932
rect 56045 13923 56103 13929
rect 54956 13892 55628 13920
rect 51905 13855 51963 13861
rect 50724 13824 51856 13852
rect 50525 13815 50583 13821
rect 47268 13756 47992 13784
rect 51828 13784 51856 13824
rect 51905 13821 51917 13855
rect 51951 13821 51963 13855
rect 51905 13815 51963 13821
rect 51997 13855 52055 13861
rect 51997 13821 52009 13855
rect 52043 13852 52055 13855
rect 52546 13852 52552 13864
rect 52043 13824 52552 13852
rect 52043 13821 52055 13824
rect 51997 13815 52055 13821
rect 52546 13812 52552 13824
rect 52604 13812 52610 13864
rect 54018 13852 54024 13864
rect 53979 13824 54024 13852
rect 54018 13812 54024 13824
rect 54076 13812 54082 13864
rect 54570 13812 54576 13864
rect 54628 13852 54634 13864
rect 54956 13852 54984 13892
rect 55490 13852 55496 13864
rect 54628 13824 54984 13852
rect 55451 13824 55496 13852
rect 54628 13812 54634 13824
rect 55490 13812 55496 13824
rect 55548 13812 55554 13864
rect 55600 13861 55628 13892
rect 56045 13889 56057 13923
rect 56091 13920 56103 13923
rect 57330 13920 57336 13932
rect 56091 13892 57336 13920
rect 56091 13889 56103 13892
rect 56045 13883 56103 13889
rect 57330 13880 57336 13892
rect 57388 13880 57394 13932
rect 55585 13855 55643 13861
rect 55585 13821 55597 13855
rect 55631 13821 55643 13855
rect 55585 13815 55643 13821
rect 53558 13784 53564 13796
rect 51828 13756 53564 13784
rect 47268 13744 47274 13756
rect 53558 13744 53564 13756
rect 53616 13744 53622 13796
rect 53926 13784 53932 13796
rect 53887 13756 53932 13784
rect 53926 13744 53932 13756
rect 53984 13744 53990 13796
rect 46198 13716 46204 13728
rect 39224 13688 46204 13716
rect 38528 13676 38534 13688
rect 46198 13676 46204 13688
rect 46256 13676 46262 13728
rect 48130 13676 48136 13728
rect 48188 13716 48194 13728
rect 49145 13719 49203 13725
rect 49145 13716 49157 13719
rect 48188 13688 49157 13716
rect 48188 13676 48194 13688
rect 49145 13685 49157 13688
rect 49191 13716 49203 13719
rect 50062 13716 50068 13728
rect 49191 13688 50068 13716
rect 49191 13685 49203 13688
rect 49145 13679 49203 13685
rect 50062 13676 50068 13688
rect 50120 13676 50126 13728
rect 1104 13626 62192 13648
rect 1104 13574 21344 13626
rect 21396 13574 21408 13626
rect 21460 13574 21472 13626
rect 21524 13574 21536 13626
rect 21588 13574 41707 13626
rect 41759 13574 41771 13626
rect 41823 13574 41835 13626
rect 41887 13574 41899 13626
rect 41951 13574 62192 13626
rect 1104 13552 62192 13574
rect 4062 13472 4068 13524
rect 4120 13512 4126 13524
rect 18874 13512 18880 13524
rect 4120 13484 18880 13512
rect 4120 13472 4126 13484
rect 18874 13472 18880 13484
rect 18932 13472 18938 13524
rect 19058 13472 19064 13524
rect 19116 13512 19122 13524
rect 22646 13512 22652 13524
rect 19116 13484 22652 13512
rect 19116 13472 19122 13484
rect 22646 13472 22652 13484
rect 22704 13472 22710 13524
rect 24394 13512 24400 13524
rect 22756 13484 24400 13512
rect 5350 13444 5356 13456
rect 5311 13416 5356 13444
rect 5350 13404 5356 13416
rect 5408 13404 5414 13456
rect 10410 13444 10416 13456
rect 10371 13416 10416 13444
rect 10410 13404 10416 13416
rect 10468 13404 10474 13456
rect 11425 13447 11483 13453
rect 11425 13413 11437 13447
rect 11471 13444 11483 13447
rect 15378 13444 15384 13456
rect 11471 13416 15384 13444
rect 11471 13413 11483 13416
rect 11425 13407 11483 13413
rect 15378 13404 15384 13416
rect 15436 13404 15442 13456
rect 17126 13444 17132 13456
rect 17087 13416 17132 13444
rect 17126 13404 17132 13416
rect 17184 13404 17190 13456
rect 18782 13404 18788 13456
rect 18840 13444 18846 13456
rect 18969 13447 19027 13453
rect 18969 13444 18981 13447
rect 18840 13416 18981 13444
rect 18840 13404 18846 13416
rect 18969 13413 18981 13416
rect 19015 13413 19027 13447
rect 20898 13444 20904 13456
rect 20859 13416 20904 13444
rect 18969 13407 19027 13413
rect 20898 13404 20904 13416
rect 20956 13404 20962 13456
rect 22756 13444 22784 13484
rect 24394 13472 24400 13484
rect 24452 13472 24458 13524
rect 25501 13515 25559 13521
rect 25501 13481 25513 13515
rect 25547 13512 25559 13515
rect 26786 13512 26792 13524
rect 25547 13484 26792 13512
rect 25547 13481 25559 13484
rect 25501 13475 25559 13481
rect 26786 13472 26792 13484
rect 26844 13472 26850 13524
rect 26878 13472 26884 13524
rect 26936 13512 26942 13524
rect 42886 13512 42892 13524
rect 26936 13484 37872 13512
rect 42847 13484 42892 13512
rect 26936 13472 26942 13484
rect 26513 13447 26571 13453
rect 26513 13444 26525 13447
rect 21560 13416 22784 13444
rect 23124 13416 26525 13444
rect 5258 13376 5264 13388
rect 5219 13348 5264 13376
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 5442 13336 5448 13388
rect 5500 13376 5506 13388
rect 9766 13376 9772 13388
rect 5500 13348 5545 13376
rect 9727 13348 9772 13376
rect 5500 13336 5506 13348
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 10134 13376 10140 13388
rect 10095 13348 10140 13376
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 12069 13379 12127 13385
rect 12069 13345 12081 13379
rect 12115 13345 12127 13379
rect 12069 13339 12127 13345
rect 11054 13268 11060 13320
rect 11112 13308 11118 13320
rect 11974 13308 11980 13320
rect 11112 13280 11980 13308
rect 11112 13268 11118 13280
rect 11974 13268 11980 13280
rect 12032 13268 12038 13320
rect 12084 13240 12112 13339
rect 12250 13336 12256 13388
rect 12308 13376 12314 13388
rect 12437 13379 12495 13385
rect 12437 13376 12449 13379
rect 12308 13348 12449 13376
rect 12308 13336 12314 13348
rect 12437 13345 12449 13348
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 13541 13379 13599 13385
rect 13541 13345 13553 13379
rect 13587 13376 13599 13379
rect 14642 13376 14648 13388
rect 13587 13348 14648 13376
rect 13587 13345 13599 13348
rect 13541 13339 13599 13345
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 15286 13376 15292 13388
rect 15247 13348 15292 13376
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 17034 13336 17040 13388
rect 17092 13376 17098 13388
rect 17589 13379 17647 13385
rect 17589 13376 17601 13379
rect 17092 13348 17601 13376
rect 17092 13336 17098 13348
rect 17589 13345 17601 13348
rect 17635 13345 17647 13379
rect 17954 13376 17960 13388
rect 17915 13348 17960 13376
rect 17589 13339 17647 13345
rect 17954 13336 17960 13348
rect 18012 13336 18018 13388
rect 19429 13379 19487 13385
rect 19429 13345 19441 13379
rect 19475 13376 19487 13379
rect 19518 13376 19524 13388
rect 19475 13348 19524 13376
rect 19475 13345 19487 13348
rect 19429 13339 19487 13345
rect 19518 13336 19524 13348
rect 19576 13336 19582 13388
rect 19794 13376 19800 13388
rect 19755 13348 19800 13376
rect 19794 13336 19800 13348
rect 19852 13336 19858 13388
rect 21174 13336 21180 13388
rect 21232 13376 21238 13388
rect 21560 13385 21588 13416
rect 21361 13379 21419 13385
rect 21361 13376 21373 13379
rect 21232 13348 21373 13376
rect 21232 13336 21238 13348
rect 21361 13345 21373 13348
rect 21407 13345 21419 13379
rect 21361 13339 21419 13345
rect 21545 13379 21603 13385
rect 21545 13345 21557 13379
rect 21591 13345 21603 13379
rect 21726 13376 21732 13388
rect 21687 13348 21732 13376
rect 21545 13339 21603 13345
rect 12342 13268 12348 13320
rect 12400 13308 12406 13320
rect 12529 13311 12587 13317
rect 12529 13308 12541 13311
rect 12400 13280 12541 13308
rect 12400 13268 12406 13280
rect 12529 13277 12541 13280
rect 12575 13308 12587 13311
rect 13262 13308 13268 13320
rect 12575 13280 13268 13308
rect 12575 13277 12587 13280
rect 12529 13271 12587 13277
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 13446 13308 13452 13320
rect 13407 13280 13452 13308
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 18049 13311 18107 13317
rect 13556 13280 15608 13308
rect 12894 13240 12900 13252
rect 12084 13212 12900 13240
rect 12894 13200 12900 13212
rect 12952 13200 12958 13252
rect 13556 13240 13584 13280
rect 13004 13212 13584 13240
rect 5534 13132 5540 13184
rect 5592 13172 5598 13184
rect 5629 13175 5687 13181
rect 5629 13172 5641 13175
rect 5592 13144 5641 13172
rect 5592 13132 5598 13144
rect 5629 13141 5641 13144
rect 5675 13141 5687 13175
rect 5629 13135 5687 13141
rect 10134 13132 10140 13184
rect 10192 13172 10198 13184
rect 13004 13172 13032 13212
rect 13630 13200 13636 13252
rect 13688 13240 13694 13252
rect 15473 13243 15531 13249
rect 15473 13240 15485 13243
rect 13688 13212 15485 13240
rect 13688 13200 13694 13212
rect 15473 13209 15485 13212
rect 15519 13209 15531 13243
rect 15473 13203 15531 13209
rect 10192 13144 13032 13172
rect 10192 13132 10198 13144
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 13725 13175 13783 13181
rect 13725 13172 13737 13175
rect 13136 13144 13737 13172
rect 13136 13132 13142 13144
rect 13725 13141 13737 13144
rect 13771 13141 13783 13175
rect 15580 13172 15608 13280
rect 18049 13277 18061 13311
rect 18095 13308 18107 13311
rect 19889 13311 19947 13317
rect 19889 13308 19901 13311
rect 18095 13280 19901 13308
rect 18095 13277 18107 13280
rect 18049 13271 18107 13277
rect 19889 13277 19901 13280
rect 19935 13308 19947 13311
rect 21560 13308 21588 13339
rect 21726 13336 21732 13348
rect 21784 13376 21790 13388
rect 22741 13379 22799 13385
rect 22741 13376 22753 13379
rect 21784 13348 22753 13376
rect 21784 13336 21790 13348
rect 22741 13345 22753 13348
rect 22787 13345 22799 13379
rect 22741 13339 22799 13345
rect 22833 13379 22891 13385
rect 22833 13345 22845 13379
rect 22879 13376 22891 13379
rect 23014 13376 23020 13388
rect 22879 13348 23020 13376
rect 22879 13345 22891 13348
rect 22833 13339 22891 13345
rect 23014 13336 23020 13348
rect 23072 13336 23078 13388
rect 23124 13308 23152 13416
rect 26513 13413 26525 13416
rect 26559 13413 26571 13447
rect 26513 13407 26571 13413
rect 28353 13447 28411 13453
rect 28353 13413 28365 13447
rect 28399 13444 28411 13447
rect 28399 13416 31984 13444
rect 28399 13413 28411 13416
rect 28353 13407 28411 13413
rect 24121 13379 24179 13385
rect 24121 13345 24133 13379
rect 24167 13376 24179 13379
rect 24210 13376 24216 13388
rect 24167 13348 24216 13376
rect 24167 13345 24179 13348
rect 24121 13339 24179 13345
rect 24210 13336 24216 13348
rect 24268 13336 24274 13388
rect 25222 13336 25228 13388
rect 25280 13376 25286 13388
rect 25317 13379 25375 13385
rect 25317 13376 25329 13379
rect 25280 13348 25329 13376
rect 25280 13336 25286 13348
rect 25317 13345 25329 13348
rect 25363 13345 25375 13379
rect 27062 13376 27068 13388
rect 27023 13348 27068 13376
rect 25317 13339 25375 13345
rect 27062 13336 27068 13348
rect 27120 13336 27126 13388
rect 27338 13376 27344 13388
rect 27299 13348 27344 13376
rect 27338 13336 27344 13348
rect 27396 13336 27402 13388
rect 27982 13336 27988 13388
rect 28040 13376 28046 13388
rect 28537 13379 28595 13385
rect 28537 13376 28549 13379
rect 28040 13348 28549 13376
rect 28040 13336 28046 13348
rect 28537 13345 28549 13348
rect 28583 13345 28595 13379
rect 30374 13376 30380 13388
rect 30335 13348 30380 13376
rect 28537 13339 28595 13345
rect 30374 13336 30380 13348
rect 30432 13336 30438 13388
rect 30561 13379 30619 13385
rect 30561 13345 30573 13379
rect 30607 13345 30619 13379
rect 30742 13376 30748 13388
rect 30703 13348 30748 13376
rect 30561 13339 30619 13345
rect 19935 13280 21588 13308
rect 21836 13280 23152 13308
rect 27525 13311 27583 13317
rect 19935 13277 19947 13280
rect 19889 13271 19947 13277
rect 17218 13200 17224 13252
rect 17276 13240 17282 13252
rect 21836 13240 21864 13280
rect 27525 13277 27537 13311
rect 27571 13308 27583 13311
rect 28258 13308 28264 13320
rect 27571 13280 28264 13308
rect 27571 13277 27583 13280
rect 27525 13271 27583 13277
rect 28258 13268 28264 13280
rect 28316 13268 28322 13320
rect 28442 13268 28448 13320
rect 28500 13308 28506 13320
rect 30576 13308 30604 13339
rect 30742 13336 30748 13348
rect 30800 13336 30806 13388
rect 28500 13280 30604 13308
rect 31956 13308 31984 13416
rect 32030 13404 32036 13456
rect 32088 13444 32094 13456
rect 32309 13447 32367 13453
rect 32309 13444 32321 13447
rect 32088 13416 32321 13444
rect 32088 13404 32094 13416
rect 32309 13413 32321 13416
rect 32355 13413 32367 13447
rect 32309 13407 32367 13413
rect 33873 13447 33931 13453
rect 33873 13413 33885 13447
rect 33919 13444 33931 13447
rect 34882 13444 34888 13456
rect 33919 13416 34888 13444
rect 33919 13413 33931 13416
rect 33873 13407 33931 13413
rect 34882 13404 34888 13416
rect 34940 13404 34946 13456
rect 36633 13447 36691 13453
rect 36633 13413 36645 13447
rect 36679 13444 36691 13447
rect 36814 13444 36820 13456
rect 36679 13416 36820 13444
rect 36679 13413 36691 13416
rect 36633 13407 36691 13413
rect 36814 13404 36820 13416
rect 36872 13404 36878 13456
rect 37734 13444 37740 13456
rect 37695 13416 37740 13444
rect 37734 13404 37740 13416
rect 37792 13404 37798 13456
rect 37844 13444 37872 13484
rect 42886 13472 42892 13484
rect 42944 13472 42950 13524
rect 53926 13472 53932 13524
rect 53984 13512 53990 13524
rect 54941 13515 54999 13521
rect 54941 13512 54953 13515
rect 53984 13484 54953 13512
rect 53984 13472 53990 13484
rect 54941 13481 54953 13484
rect 54987 13481 54999 13515
rect 54941 13475 54999 13481
rect 41322 13444 41328 13456
rect 37844 13416 41328 13444
rect 41322 13404 41328 13416
rect 41380 13404 41386 13456
rect 41509 13447 41567 13453
rect 41509 13413 41521 13447
rect 41555 13444 41567 13447
rect 42058 13444 42064 13456
rect 41555 13416 42064 13444
rect 41555 13413 41567 13416
rect 41509 13407 41567 13413
rect 42058 13404 42064 13416
rect 42116 13404 42122 13456
rect 44545 13447 44603 13453
rect 44545 13413 44557 13447
rect 44591 13444 44603 13447
rect 45278 13444 45284 13456
rect 44591 13416 45284 13444
rect 44591 13413 44603 13416
rect 44545 13407 44603 13413
rect 45278 13404 45284 13416
rect 45336 13404 45342 13456
rect 48961 13447 49019 13453
rect 48961 13413 48973 13447
rect 49007 13444 49019 13447
rect 49234 13444 49240 13456
rect 49007 13416 49240 13444
rect 49007 13413 49019 13416
rect 48961 13407 49019 13413
rect 49234 13404 49240 13416
rect 49292 13404 49298 13456
rect 52457 13447 52515 13453
rect 52457 13413 52469 13447
rect 52503 13444 52515 13447
rect 53006 13444 53012 13456
rect 52503 13416 53012 13444
rect 52503 13413 52515 13416
rect 52457 13407 52515 13413
rect 53006 13404 53012 13416
rect 53064 13404 53070 13456
rect 54662 13444 54668 13456
rect 54623 13416 54668 13444
rect 54662 13404 54668 13416
rect 54720 13404 54726 13456
rect 32398 13376 32404 13388
rect 32359 13348 32404 13376
rect 32398 13336 32404 13348
rect 32456 13336 32462 13388
rect 33965 13379 34023 13385
rect 33965 13345 33977 13379
rect 34011 13345 34023 13379
rect 33965 13339 34023 13345
rect 33870 13308 33876 13320
rect 31956 13280 33876 13308
rect 28500 13268 28506 13280
rect 33870 13268 33876 13280
rect 33928 13268 33934 13320
rect 26234 13240 26240 13252
rect 17276 13212 21864 13240
rect 22756 13212 26240 13240
rect 17276 13200 17282 13212
rect 22756 13172 22784 13212
rect 26234 13200 26240 13212
rect 26292 13200 26298 13252
rect 30098 13240 30104 13252
rect 28552 13212 30104 13240
rect 15580 13144 22784 13172
rect 13725 13135 13783 13141
rect 22830 13132 22836 13184
rect 22888 13172 22894 13184
rect 23017 13175 23075 13181
rect 23017 13172 23029 13175
rect 22888 13144 23029 13172
rect 22888 13132 22894 13144
rect 23017 13141 23029 13144
rect 23063 13141 23075 13175
rect 24302 13172 24308 13184
rect 24263 13144 24308 13172
rect 23017 13135 23075 13141
rect 24302 13132 24308 13144
rect 24360 13132 24366 13184
rect 25774 13132 25780 13184
rect 25832 13172 25838 13184
rect 28552 13172 28580 13212
rect 30098 13200 30104 13212
rect 30156 13200 30162 13252
rect 30193 13243 30251 13249
rect 30193 13209 30205 13243
rect 30239 13240 30251 13243
rect 30466 13240 30472 13252
rect 30239 13212 30472 13240
rect 30239 13209 30251 13212
rect 30193 13203 30251 13209
rect 30466 13200 30472 13212
rect 30524 13200 30530 13252
rect 31110 13200 31116 13252
rect 31168 13240 31174 13252
rect 33980 13240 34008 13339
rect 35158 13336 35164 13388
rect 35216 13376 35222 13388
rect 36170 13376 36176 13388
rect 35216 13348 36176 13376
rect 35216 13336 35222 13348
rect 36170 13336 36176 13348
rect 36228 13336 36234 13388
rect 38378 13376 38384 13388
rect 38339 13348 38384 13376
rect 38378 13336 38384 13348
rect 38436 13336 38442 13388
rect 38470 13336 38476 13388
rect 38528 13376 38534 13388
rect 38749 13379 38807 13385
rect 38528 13348 38573 13376
rect 38528 13336 38534 13348
rect 38749 13345 38761 13379
rect 38795 13345 38807 13379
rect 38749 13339 38807 13345
rect 38933 13379 38991 13385
rect 38933 13345 38945 13379
rect 38979 13376 38991 13379
rect 39390 13376 39396 13388
rect 38979 13348 39396 13376
rect 38979 13345 38991 13348
rect 38933 13339 38991 13345
rect 35066 13268 35072 13320
rect 35124 13308 35130 13320
rect 36081 13311 36139 13317
rect 36081 13308 36093 13311
rect 35124 13280 36093 13308
rect 35124 13268 35130 13280
rect 36081 13277 36093 13280
rect 36127 13277 36139 13311
rect 36081 13271 36139 13277
rect 36354 13240 36360 13252
rect 31168 13212 32628 13240
rect 33980 13212 36360 13240
rect 31168 13200 31174 13212
rect 25832 13144 28580 13172
rect 28629 13175 28687 13181
rect 25832 13132 25838 13144
rect 28629 13141 28641 13175
rect 28675 13172 28687 13175
rect 28718 13172 28724 13184
rect 28675 13144 28724 13172
rect 28675 13141 28687 13144
rect 28629 13135 28687 13141
rect 28718 13132 28724 13144
rect 28776 13132 28782 13184
rect 30282 13132 30288 13184
rect 30340 13172 30346 13184
rect 30926 13172 30932 13184
rect 30340 13144 30932 13172
rect 30340 13132 30346 13144
rect 30926 13132 30932 13144
rect 30984 13172 30990 13184
rect 32600 13181 32628 13212
rect 36354 13200 36360 13212
rect 36412 13200 36418 13252
rect 38764 13240 38792 13339
rect 39390 13336 39396 13348
rect 39448 13336 39454 13388
rect 41598 13336 41604 13388
rect 41656 13376 41662 13388
rect 41693 13379 41751 13385
rect 41693 13376 41705 13379
rect 41656 13348 41705 13376
rect 41656 13336 41662 13348
rect 41693 13345 41705 13348
rect 41739 13345 41751 13379
rect 43070 13376 43076 13388
rect 43031 13348 43076 13376
rect 41693 13339 41751 13345
rect 41708 13308 41736 13339
rect 43070 13336 43076 13348
rect 43128 13336 43134 13388
rect 43162 13336 43168 13388
rect 43220 13376 43226 13388
rect 45189 13379 45247 13385
rect 45189 13376 45201 13379
rect 43220 13348 45201 13376
rect 43220 13336 43226 13348
rect 45189 13345 45201 13348
rect 45235 13345 45247 13379
rect 45189 13339 45247 13345
rect 45557 13379 45615 13385
rect 45557 13345 45569 13379
rect 45603 13376 45615 13379
rect 45738 13376 45744 13388
rect 45603 13348 45744 13376
rect 45603 13345 45615 13348
rect 45557 13339 45615 13345
rect 45738 13336 45744 13348
rect 45796 13336 45802 13388
rect 46106 13336 46112 13388
rect 46164 13376 46170 13388
rect 46753 13379 46811 13385
rect 46753 13376 46765 13379
rect 46164 13348 46765 13376
rect 46164 13336 46170 13348
rect 46753 13345 46765 13348
rect 46799 13345 46811 13379
rect 46753 13339 46811 13345
rect 47118 13336 47124 13388
rect 47176 13376 47182 13388
rect 47489 13379 47547 13385
rect 47489 13376 47501 13379
rect 47176 13348 47501 13376
rect 47176 13336 47182 13348
rect 47489 13345 47501 13348
rect 47535 13345 47547 13379
rect 47489 13339 47547 13345
rect 47578 13336 47584 13388
rect 47636 13376 47642 13388
rect 47857 13379 47915 13385
rect 47857 13376 47869 13379
rect 47636 13348 47869 13376
rect 47636 13336 47642 13348
rect 47857 13345 47869 13348
rect 47903 13345 47915 13379
rect 47857 13339 47915 13345
rect 48041 13379 48099 13385
rect 48041 13345 48053 13379
rect 48087 13376 48099 13379
rect 48130 13376 48136 13388
rect 48087 13348 48136 13376
rect 48087 13345 48099 13348
rect 48041 13339 48099 13345
rect 44358 13308 44364 13320
rect 41708 13280 44364 13308
rect 44358 13268 44364 13280
rect 44416 13268 44422 13320
rect 44726 13268 44732 13320
rect 44784 13308 44790 13320
rect 45097 13311 45155 13317
rect 45097 13308 45109 13311
rect 44784 13280 45109 13308
rect 44784 13268 44790 13280
rect 45097 13277 45109 13280
rect 45143 13277 45155 13311
rect 45646 13308 45652 13320
rect 45559 13280 45652 13308
rect 45097 13271 45155 13277
rect 45646 13268 45652 13280
rect 45704 13308 45710 13320
rect 45830 13308 45836 13320
rect 45704 13280 45836 13308
rect 45704 13268 45710 13280
rect 45830 13268 45836 13280
rect 45888 13308 45894 13320
rect 45888 13280 47348 13308
rect 45888 13268 45894 13280
rect 46474 13240 46480 13252
rect 38764 13212 46480 13240
rect 46474 13200 46480 13212
rect 46532 13200 46538 13252
rect 46934 13240 46940 13252
rect 46895 13212 46940 13240
rect 46934 13200 46940 13212
rect 46992 13200 46998 13252
rect 47320 13240 47348 13280
rect 47394 13268 47400 13320
rect 47452 13308 47458 13320
rect 47452 13280 47497 13308
rect 47452 13268 47458 13280
rect 48056 13240 48084 13339
rect 48130 13336 48136 13348
rect 48188 13336 48194 13388
rect 49602 13376 49608 13388
rect 49563 13348 49608 13376
rect 49602 13336 49608 13348
rect 49660 13336 49666 13388
rect 49970 13376 49976 13388
rect 49931 13348 49976 13376
rect 49970 13336 49976 13348
rect 50028 13336 50034 13388
rect 51166 13376 51172 13388
rect 51127 13348 51172 13376
rect 51166 13336 51172 13348
rect 51224 13336 51230 13388
rect 53098 13376 53104 13388
rect 53059 13348 53104 13376
rect 53098 13336 53104 13348
rect 53156 13336 53162 13388
rect 53374 13336 53380 13388
rect 53432 13385 53438 13388
rect 53432 13379 53493 13385
rect 53432 13345 53447 13379
rect 53481 13345 53493 13379
rect 53432 13339 53493 13345
rect 54849 13379 54907 13385
rect 54849 13345 54861 13379
rect 54895 13376 54907 13379
rect 56502 13376 56508 13388
rect 54895 13348 56508 13376
rect 54895 13345 54907 13348
rect 54849 13339 54907 13345
rect 53432 13336 53438 13339
rect 56502 13336 56508 13348
rect 56560 13336 56566 13388
rect 48222 13268 48228 13320
rect 48280 13308 48286 13320
rect 49513 13311 49571 13317
rect 49513 13308 49525 13311
rect 48280 13280 49525 13308
rect 48280 13268 48286 13280
rect 49513 13277 49525 13280
rect 49559 13277 49571 13311
rect 50062 13308 50068 13320
rect 50023 13280 50068 13308
rect 49513 13271 49571 13277
rect 50062 13268 50068 13280
rect 50120 13268 50126 13320
rect 50614 13268 50620 13320
rect 50672 13308 50678 13320
rect 51077 13311 51135 13317
rect 51077 13308 51089 13311
rect 50672 13280 51089 13308
rect 50672 13268 50678 13280
rect 51077 13277 51089 13280
rect 51123 13277 51135 13311
rect 51626 13308 51632 13320
rect 51587 13280 51632 13308
rect 51077 13271 51135 13277
rect 51626 13268 51632 13280
rect 51684 13268 51690 13320
rect 53190 13308 53196 13320
rect 53151 13280 53196 13308
rect 53190 13268 53196 13280
rect 53248 13268 53254 13320
rect 53558 13308 53564 13320
rect 53519 13280 53564 13308
rect 53558 13268 53564 13280
rect 53616 13268 53622 13320
rect 47320 13212 48084 13240
rect 32125 13175 32183 13181
rect 32125 13172 32137 13175
rect 30984 13144 32137 13172
rect 30984 13132 30990 13144
rect 32125 13141 32137 13144
rect 32171 13141 32183 13175
rect 32125 13135 32183 13141
rect 32585 13175 32643 13181
rect 32585 13141 32597 13175
rect 32631 13141 32643 13175
rect 33686 13172 33692 13184
rect 33647 13144 33692 13172
rect 32585 13135 32643 13141
rect 33686 13132 33692 13144
rect 33744 13132 33750 13184
rect 33778 13132 33784 13184
rect 33836 13172 33842 13184
rect 34149 13175 34207 13181
rect 34149 13172 34161 13175
rect 33836 13144 34161 13172
rect 33836 13132 33842 13144
rect 34149 13141 34161 13144
rect 34195 13141 34207 13175
rect 34149 13135 34207 13141
rect 34238 13132 34244 13184
rect 34296 13172 34302 13184
rect 40494 13172 40500 13184
rect 34296 13144 40500 13172
rect 34296 13132 34302 13144
rect 40494 13132 40500 13144
rect 40552 13132 40558 13184
rect 41414 13132 41420 13184
rect 41472 13172 41478 13184
rect 41785 13175 41843 13181
rect 41785 13172 41797 13175
rect 41472 13144 41797 13172
rect 41472 13132 41478 13144
rect 41785 13141 41797 13144
rect 41831 13141 41843 13175
rect 41785 13135 41843 13141
rect 45922 13132 45928 13184
rect 45980 13172 45986 13184
rect 46569 13175 46627 13181
rect 46569 13172 46581 13175
rect 45980 13144 46581 13172
rect 45980 13132 45986 13144
rect 46569 13141 46581 13144
rect 46615 13172 46627 13175
rect 46658 13172 46664 13184
rect 46615 13144 46664 13172
rect 46615 13141 46627 13144
rect 46569 13135 46627 13141
rect 46658 13132 46664 13144
rect 46716 13132 46722 13184
rect 1104 13082 62192 13104
rect 1104 13030 11163 13082
rect 11215 13030 11227 13082
rect 11279 13030 11291 13082
rect 11343 13030 11355 13082
rect 11407 13030 31526 13082
rect 31578 13030 31590 13082
rect 31642 13030 31654 13082
rect 31706 13030 31718 13082
rect 31770 13030 51888 13082
rect 51940 13030 51952 13082
rect 52004 13030 52016 13082
rect 52068 13030 52080 13082
rect 52132 13030 62192 13082
rect 1104 13008 62192 13030
rect 4801 12971 4859 12977
rect 4801 12937 4813 12971
rect 4847 12968 4859 12971
rect 5442 12968 5448 12980
rect 4847 12940 5448 12968
rect 4847 12937 4859 12940
rect 4801 12931 4859 12937
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 10413 12971 10471 12977
rect 5552 12940 9076 12968
rect 3050 12860 3056 12912
rect 3108 12900 3114 12912
rect 5552 12900 5580 12940
rect 8938 12900 8944 12912
rect 3108 12872 5580 12900
rect 5736 12872 8944 12900
rect 3108 12860 3114 12872
rect 5353 12767 5411 12773
rect 5353 12733 5365 12767
rect 5399 12733 5411 12767
rect 5353 12727 5411 12733
rect 5445 12767 5503 12773
rect 5445 12733 5457 12767
rect 5491 12764 5503 12767
rect 5626 12764 5632 12776
rect 5491 12736 5632 12764
rect 5491 12733 5503 12736
rect 5445 12727 5503 12733
rect 5368 12696 5396 12727
rect 5626 12724 5632 12736
rect 5684 12724 5690 12776
rect 5736 12773 5764 12872
rect 8938 12860 8944 12872
rect 8996 12860 9002 12912
rect 9048 12900 9076 12940
rect 10413 12937 10425 12971
rect 10459 12968 10471 12971
rect 12618 12968 12624 12980
rect 10459 12940 12624 12968
rect 10459 12937 10471 12940
rect 10413 12931 10471 12937
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 17218 12968 17224 12980
rect 12820 12940 17224 12968
rect 12820 12900 12848 12940
rect 17218 12928 17224 12940
rect 17276 12928 17282 12980
rect 18138 12928 18144 12980
rect 18196 12968 18202 12980
rect 18233 12971 18291 12977
rect 18233 12968 18245 12971
rect 18196 12940 18245 12968
rect 18196 12928 18202 12940
rect 18233 12937 18245 12940
rect 18279 12968 18291 12971
rect 20346 12968 20352 12980
rect 18279 12940 20352 12968
rect 18279 12937 18291 12940
rect 18233 12931 18291 12937
rect 20346 12928 20352 12940
rect 20404 12928 20410 12980
rect 22281 12971 22339 12977
rect 22281 12968 22293 12971
rect 20548 12940 22293 12968
rect 9048 12872 12848 12900
rect 12912 12872 16620 12900
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 7282 12832 7288 12844
rect 6871 12804 7288 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12832 7435 12835
rect 8294 12832 8300 12844
rect 7423 12804 8300 12832
rect 7423 12801 7435 12804
rect 7377 12795 7435 12801
rect 8294 12792 8300 12804
rect 8352 12792 8358 12844
rect 12912 12832 12940 12872
rect 8404 12804 12940 12832
rect 12989 12835 13047 12841
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12733 5779 12767
rect 5721 12727 5779 12733
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12764 5963 12767
rect 6454 12764 6460 12776
rect 5951 12736 6460 12764
rect 5951 12733 5963 12736
rect 5905 12727 5963 12733
rect 6454 12724 6460 12736
rect 6512 12724 6518 12776
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12764 6975 12767
rect 7466 12764 7472 12776
rect 6963 12736 7472 12764
rect 6963 12733 6975 12736
rect 6917 12727 6975 12733
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 7006 12696 7012 12708
rect 5368 12668 7012 12696
rect 7006 12656 7012 12668
rect 7064 12656 7070 12708
rect 6546 12588 6552 12640
rect 6604 12628 6610 12640
rect 8404 12628 8432 12804
rect 12989 12801 13001 12835
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 9214 12764 9220 12776
rect 9175 12736 9220 12764
rect 9214 12724 9220 12736
rect 9272 12724 9278 12776
rect 9306 12724 9312 12776
rect 9364 12764 9370 12776
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 9364 12736 10977 12764
rect 9364 12724 9370 12736
rect 10965 12733 10977 12736
rect 11011 12733 11023 12767
rect 10965 12727 11023 12733
rect 11054 12724 11060 12776
rect 11112 12764 11118 12776
rect 11333 12767 11391 12773
rect 11112 12736 11205 12764
rect 11112 12724 11118 12736
rect 11333 12733 11345 12767
rect 11379 12733 11391 12767
rect 11514 12764 11520 12776
rect 11475 12736 11520 12764
rect 11333 12727 11391 12733
rect 11072 12696 11100 12724
rect 11238 12696 11244 12708
rect 10980 12668 11244 12696
rect 6604 12600 8432 12628
rect 9401 12631 9459 12637
rect 6604 12588 6610 12600
rect 9401 12597 9413 12631
rect 9447 12628 9459 12631
rect 10980 12628 11008 12668
rect 11238 12656 11244 12668
rect 11296 12656 11302 12708
rect 9447 12600 11008 12628
rect 11348 12628 11376 12727
rect 11514 12724 11520 12736
rect 11572 12724 11578 12776
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 13004 12764 13032 12795
rect 13262 12792 13268 12844
rect 13320 12832 13326 12844
rect 13541 12835 13599 12841
rect 13541 12832 13553 12835
rect 13320 12804 13553 12832
rect 13320 12792 13326 12804
rect 13541 12801 13553 12804
rect 13587 12801 13599 12835
rect 13541 12795 13599 12801
rect 12032 12736 13032 12764
rect 12032 12724 12038 12736
rect 13078 12724 13084 12776
rect 13136 12764 13142 12776
rect 13136 12736 13181 12764
rect 13136 12724 13142 12736
rect 13354 12724 13360 12776
rect 13412 12764 13418 12776
rect 13449 12767 13507 12773
rect 13449 12764 13461 12767
rect 13412 12736 13461 12764
rect 13412 12724 13418 12736
rect 13449 12733 13461 12736
rect 13495 12733 13507 12767
rect 13449 12727 13507 12733
rect 13998 12724 14004 12776
rect 14056 12764 14062 12776
rect 14461 12767 14519 12773
rect 14461 12764 14473 12767
rect 14056 12736 14473 12764
rect 14056 12724 14062 12736
rect 14461 12733 14473 12736
rect 14507 12733 14519 12767
rect 15746 12764 15752 12776
rect 15707 12736 15752 12764
rect 14461 12727 14519 12733
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 16592 12773 16620 12872
rect 17586 12860 17592 12912
rect 17644 12900 17650 12912
rect 19610 12900 19616 12912
rect 17644 12872 19616 12900
rect 17644 12860 17650 12872
rect 19610 12860 19616 12872
rect 19668 12900 19674 12912
rect 20438 12900 20444 12912
rect 19668 12872 20444 12900
rect 19668 12860 19674 12872
rect 20438 12860 20444 12872
rect 20496 12860 20502 12912
rect 20548 12841 20576 12940
rect 22281 12937 22293 12940
rect 22327 12937 22339 12971
rect 22281 12931 22339 12937
rect 24302 12928 24308 12980
rect 24360 12968 24366 12980
rect 29365 12971 29423 12977
rect 29365 12968 29377 12971
rect 24360 12940 29377 12968
rect 24360 12928 24366 12940
rect 29365 12937 29377 12940
rect 29411 12937 29423 12971
rect 29365 12931 29423 12937
rect 29641 12971 29699 12977
rect 29641 12937 29653 12971
rect 29687 12968 29699 12971
rect 30834 12968 30840 12980
rect 29687 12940 30840 12968
rect 29687 12937 29699 12940
rect 29641 12931 29699 12937
rect 30834 12928 30840 12940
rect 30892 12928 30898 12980
rect 32030 12968 32036 12980
rect 31588 12940 31800 12968
rect 31991 12940 32036 12968
rect 23845 12903 23903 12909
rect 23845 12900 23857 12903
rect 23768 12872 23857 12900
rect 19797 12835 19855 12841
rect 19797 12832 19809 12835
rect 18432 12804 19809 12832
rect 16577 12767 16635 12773
rect 16577 12733 16589 12767
rect 16623 12733 16635 12767
rect 16577 12727 16635 12733
rect 16666 12724 16672 12776
rect 16724 12764 16730 12776
rect 16761 12767 16819 12773
rect 16761 12764 16773 12767
rect 16724 12736 16773 12764
rect 16724 12724 16730 12736
rect 16761 12733 16773 12736
rect 16807 12764 16819 12767
rect 17586 12764 17592 12776
rect 16807 12736 17592 12764
rect 16807 12733 16819 12736
rect 16761 12727 16819 12733
rect 17586 12724 17592 12736
rect 17644 12724 17650 12776
rect 18432 12773 18460 12804
rect 19797 12801 19809 12804
rect 19843 12801 19855 12835
rect 19797 12795 19855 12801
rect 20533 12835 20591 12841
rect 20533 12801 20545 12835
rect 20579 12801 20591 12835
rect 20533 12795 20591 12801
rect 20622 12792 20628 12844
rect 20680 12832 20686 12844
rect 21821 12835 21879 12841
rect 21821 12832 21833 12835
rect 20680 12804 21833 12832
rect 20680 12792 20686 12804
rect 21821 12801 21833 12804
rect 21867 12832 21879 12835
rect 23768 12832 23796 12872
rect 23845 12869 23857 12872
rect 23891 12900 23903 12903
rect 25774 12900 25780 12912
rect 23891 12872 25780 12900
rect 23891 12869 23903 12872
rect 23845 12863 23903 12869
rect 25774 12860 25780 12872
rect 25832 12860 25838 12912
rect 25869 12903 25927 12909
rect 25869 12869 25881 12903
rect 25915 12900 25927 12903
rect 26142 12900 26148 12912
rect 25915 12872 26148 12900
rect 25915 12869 25927 12872
rect 25869 12863 25927 12869
rect 26142 12860 26148 12872
rect 26200 12860 26206 12912
rect 26234 12860 26240 12912
rect 26292 12900 26298 12912
rect 31588 12900 31616 12940
rect 26292 12872 31616 12900
rect 31772 12900 31800 12940
rect 32030 12928 32036 12940
rect 32088 12928 32094 12980
rect 40586 12968 40592 12980
rect 33796 12940 40592 12968
rect 33796 12900 33824 12940
rect 40586 12928 40592 12940
rect 40644 12928 40650 12980
rect 40770 12968 40776 12980
rect 40731 12940 40776 12968
rect 40770 12928 40776 12940
rect 40828 12928 40834 12980
rect 43070 12928 43076 12980
rect 43128 12968 43134 12980
rect 45189 12971 45247 12977
rect 45189 12968 45201 12971
rect 43128 12940 45201 12968
rect 43128 12928 43134 12940
rect 45189 12937 45201 12940
rect 45235 12968 45247 12971
rect 46106 12968 46112 12980
rect 45235 12940 46112 12968
rect 45235 12937 45247 12940
rect 45189 12931 45247 12937
rect 46106 12928 46112 12940
rect 46164 12928 46170 12980
rect 46201 12971 46259 12977
rect 46201 12937 46213 12971
rect 46247 12968 46259 12971
rect 46382 12968 46388 12980
rect 46247 12940 46388 12968
rect 46247 12937 46259 12940
rect 46201 12931 46259 12937
rect 46382 12928 46388 12940
rect 46440 12928 46446 12980
rect 49602 12928 49608 12980
rect 49660 12968 49666 12980
rect 50525 12971 50583 12977
rect 50525 12968 50537 12971
rect 49660 12940 50537 12968
rect 49660 12928 49666 12940
rect 50525 12937 50537 12940
rect 50571 12937 50583 12971
rect 50525 12931 50583 12937
rect 52733 12971 52791 12977
rect 52733 12937 52745 12971
rect 52779 12968 52791 12971
rect 54018 12968 54024 12980
rect 52779 12940 54024 12968
rect 52779 12937 52791 12940
rect 52733 12931 52791 12937
rect 54018 12928 54024 12940
rect 54076 12928 54082 12980
rect 54757 12971 54815 12977
rect 54757 12937 54769 12971
rect 54803 12968 54815 12971
rect 55214 12968 55220 12980
rect 54803 12940 55220 12968
rect 54803 12937 54815 12940
rect 54757 12931 54815 12937
rect 55214 12928 55220 12940
rect 55272 12928 55278 12980
rect 47026 12900 47032 12912
rect 31772 12872 33824 12900
rect 34532 12872 43392 12900
rect 26292 12860 26298 12872
rect 26602 12832 26608 12844
rect 21867 12804 23796 12832
rect 26436 12804 26608 12832
rect 21867 12801 21879 12804
rect 21821 12795 21879 12801
rect 18417 12767 18475 12773
rect 18417 12733 18429 12767
rect 18463 12733 18475 12767
rect 18417 12727 18475 12733
rect 18509 12767 18567 12773
rect 18509 12733 18521 12767
rect 18555 12764 18567 12767
rect 20070 12764 20076 12776
rect 18555 12736 20076 12764
rect 18555 12733 18567 12736
rect 18509 12727 18567 12733
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 20254 12724 20260 12776
rect 20312 12764 20318 12776
rect 20441 12767 20499 12773
rect 20441 12764 20453 12767
rect 20312 12736 20453 12764
rect 20312 12724 20318 12736
rect 20441 12733 20453 12736
rect 20487 12733 20499 12767
rect 20806 12764 20812 12776
rect 20767 12736 20812 12764
rect 20441 12727 20499 12733
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 20901 12767 20959 12773
rect 20901 12733 20913 12767
rect 20947 12764 20959 12767
rect 20947 12736 21128 12764
rect 20947 12733 20959 12736
rect 20901 12727 20959 12733
rect 12437 12699 12495 12705
rect 12437 12665 12449 12699
rect 12483 12696 12495 12699
rect 15194 12696 15200 12708
rect 12483 12668 15200 12696
rect 12483 12665 12495 12668
rect 12437 12659 12495 12665
rect 15194 12656 15200 12668
rect 15252 12656 15258 12708
rect 17129 12699 17187 12705
rect 15488 12668 17080 12696
rect 12526 12628 12532 12640
rect 11348 12600 12532 12628
rect 9447 12597 9459 12600
rect 9401 12591 9459 12597
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 14642 12628 14648 12640
rect 14603 12600 14648 12628
rect 14642 12588 14648 12600
rect 14700 12628 14706 12640
rect 15488 12628 15516 12668
rect 14700 12600 15516 12628
rect 15565 12631 15623 12637
rect 14700 12588 14706 12600
rect 15565 12597 15577 12631
rect 15611 12628 15623 12631
rect 16574 12628 16580 12640
rect 15611 12600 16580 12628
rect 15611 12597 15623 12600
rect 15565 12591 15623 12597
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 17052 12628 17080 12668
rect 17129 12665 17141 12699
rect 17175 12696 17187 12699
rect 18782 12696 18788 12708
rect 17175 12668 18788 12696
rect 17175 12665 17187 12668
rect 17129 12659 17187 12665
rect 18782 12656 18788 12668
rect 18840 12656 18846 12708
rect 18874 12656 18880 12708
rect 18932 12696 18938 12708
rect 18969 12699 19027 12705
rect 18969 12696 18981 12699
rect 18932 12668 18981 12696
rect 18932 12656 18938 12668
rect 18969 12665 18981 12668
rect 19015 12665 19027 12699
rect 19426 12696 19432 12708
rect 18969 12659 19027 12665
rect 19260 12668 19432 12696
rect 19260 12628 19288 12668
rect 19426 12656 19432 12668
rect 19484 12656 19490 12708
rect 17052 12600 19288 12628
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 21100 12628 21128 12736
rect 22094 12724 22100 12776
rect 22152 12764 22158 12776
rect 23658 12764 23664 12776
rect 22152 12736 22197 12764
rect 23619 12736 23664 12764
rect 22152 12724 22158 12736
rect 23658 12724 23664 12736
rect 23716 12724 23722 12776
rect 23934 12724 23940 12776
rect 23992 12764 23998 12776
rect 26436 12773 26464 12804
rect 26602 12792 26608 12804
rect 26660 12792 26666 12844
rect 28442 12832 28448 12844
rect 26712 12804 28448 12832
rect 26053 12767 26111 12773
rect 26053 12764 26065 12767
rect 23992 12736 26065 12764
rect 23992 12724 23998 12736
rect 26053 12733 26065 12736
rect 26099 12733 26111 12767
rect 26053 12727 26111 12733
rect 26421 12767 26479 12773
rect 26421 12733 26433 12767
rect 26467 12733 26479 12767
rect 26421 12727 26479 12733
rect 26513 12767 26571 12773
rect 26513 12733 26525 12767
rect 26559 12764 26571 12767
rect 26712 12764 26740 12804
rect 28442 12792 28448 12804
rect 28500 12792 28506 12844
rect 29365 12835 29423 12841
rect 29365 12801 29377 12835
rect 29411 12832 29423 12835
rect 32677 12835 32735 12841
rect 29411 12804 30788 12832
rect 29411 12801 29423 12804
rect 29365 12795 29423 12801
rect 26559 12736 26740 12764
rect 26559 12733 26571 12736
rect 26513 12727 26571 12733
rect 22005 12699 22063 12705
rect 22005 12665 22017 12699
rect 22051 12696 22063 12699
rect 26326 12696 26332 12708
rect 22051 12668 26332 12696
rect 22051 12665 22063 12668
rect 22005 12659 22063 12665
rect 26326 12656 26332 12668
rect 26384 12656 26390 12708
rect 19392 12600 21128 12628
rect 19392 12588 19398 12600
rect 24394 12588 24400 12640
rect 24452 12628 24458 12640
rect 26528 12628 26556 12727
rect 26786 12724 26792 12776
rect 26844 12764 26850 12776
rect 27617 12767 27675 12773
rect 27617 12764 27629 12767
rect 26844 12736 27629 12764
rect 26844 12724 26850 12736
rect 27617 12733 27629 12736
rect 27663 12733 27675 12767
rect 27617 12727 27675 12733
rect 27706 12724 27712 12776
rect 27764 12764 27770 12776
rect 28534 12764 28540 12776
rect 27764 12736 28540 12764
rect 27764 12724 27770 12736
rect 28534 12724 28540 12736
rect 28592 12764 28598 12776
rect 29457 12767 29515 12773
rect 29457 12764 29469 12767
rect 28592 12736 29469 12764
rect 28592 12724 28598 12736
rect 29457 12733 29469 12736
rect 29503 12733 29515 12767
rect 30650 12764 30656 12776
rect 29457 12727 29515 12733
rect 29564 12736 30656 12764
rect 27433 12699 27491 12705
rect 27433 12665 27445 12699
rect 27479 12696 27491 12699
rect 29362 12696 29368 12708
rect 27479 12668 29368 12696
rect 27479 12665 27491 12668
rect 27433 12659 27491 12665
rect 29362 12656 29368 12668
rect 29420 12656 29426 12708
rect 24452 12600 26556 12628
rect 24452 12588 24458 12600
rect 27614 12588 27620 12640
rect 27672 12628 27678 12640
rect 27709 12631 27767 12637
rect 27709 12628 27721 12631
rect 27672 12600 27721 12628
rect 27672 12588 27678 12600
rect 27709 12597 27721 12600
rect 27755 12597 27767 12631
rect 27709 12591 27767 12597
rect 27890 12588 27896 12640
rect 27948 12628 27954 12640
rect 29564 12628 29592 12736
rect 30650 12724 30656 12736
rect 30708 12724 30714 12776
rect 30760 12773 30788 12804
rect 32677 12801 32689 12835
rect 32723 12832 32735 12835
rect 34422 12832 34428 12844
rect 32723 12804 34428 12832
rect 32723 12801 32735 12804
rect 32677 12795 32735 12801
rect 34422 12792 34428 12804
rect 34480 12792 34486 12844
rect 30745 12767 30803 12773
rect 30745 12733 30757 12767
rect 30791 12764 30803 12767
rect 32582 12764 32588 12776
rect 30791 12736 32444 12764
rect 32543 12736 32588 12764
rect 30791 12733 30803 12736
rect 30745 12727 30803 12733
rect 30561 12699 30619 12705
rect 30561 12665 30573 12699
rect 30607 12696 30619 12699
rect 32416 12696 32444 12736
rect 32582 12724 32588 12736
rect 32640 12724 32646 12776
rect 32950 12764 32956 12776
rect 32911 12736 32956 12764
rect 32950 12724 32956 12736
rect 33008 12724 33014 12776
rect 33045 12767 33103 12773
rect 33045 12733 33057 12767
rect 33091 12764 33103 12767
rect 34532 12764 34560 12872
rect 36633 12835 36691 12841
rect 36633 12801 36645 12835
rect 36679 12832 36691 12835
rect 38378 12832 38384 12844
rect 36679 12804 38384 12832
rect 36679 12801 36691 12804
rect 36633 12795 36691 12801
rect 38378 12792 38384 12804
rect 38436 12792 38442 12844
rect 40494 12832 40500 12844
rect 40455 12804 40500 12832
rect 40494 12792 40500 12804
rect 40552 12792 40558 12844
rect 42521 12835 42579 12841
rect 42521 12801 42533 12835
rect 42567 12832 42579 12835
rect 43162 12832 43168 12844
rect 42567 12804 43168 12832
rect 42567 12801 42579 12804
rect 42521 12795 42579 12801
rect 43162 12792 43168 12804
rect 43220 12792 43226 12844
rect 43364 12841 43392 12872
rect 46860 12872 47032 12900
rect 43349 12835 43407 12841
rect 43349 12801 43361 12835
rect 43395 12801 43407 12835
rect 43349 12795 43407 12801
rect 43901 12835 43959 12841
rect 43901 12801 43913 12835
rect 43947 12832 43959 12835
rect 45094 12832 45100 12844
rect 43947 12804 45100 12832
rect 43947 12801 43959 12804
rect 43901 12795 43959 12801
rect 45094 12792 45100 12804
rect 45152 12792 45158 12844
rect 46860 12841 46888 12872
rect 47026 12860 47032 12872
rect 47084 12900 47090 12912
rect 48222 12900 48228 12912
rect 47084 12872 48228 12900
rect 47084 12860 47090 12872
rect 48222 12860 48228 12872
rect 48280 12900 48286 12912
rect 48317 12903 48375 12909
rect 48317 12900 48329 12903
rect 48280 12872 48329 12900
rect 48280 12860 48286 12872
rect 48317 12869 48329 12872
rect 48363 12869 48375 12903
rect 48317 12863 48375 12869
rect 46845 12835 46903 12841
rect 46845 12801 46857 12835
rect 46891 12801 46903 12835
rect 47210 12832 47216 12844
rect 47171 12804 47216 12832
rect 46845 12795 46903 12801
rect 47210 12792 47216 12804
rect 47268 12792 47274 12844
rect 53190 12832 53196 12844
rect 53151 12804 53196 12832
rect 53190 12792 53196 12804
rect 53248 12792 53254 12844
rect 53558 12792 53564 12844
rect 53616 12832 53622 12844
rect 53745 12835 53803 12841
rect 53745 12832 53757 12835
rect 53616 12804 53757 12832
rect 53616 12792 53622 12804
rect 53745 12801 53757 12804
rect 53791 12801 53803 12835
rect 53745 12795 53803 12801
rect 55030 12792 55036 12844
rect 55088 12832 55094 12844
rect 55217 12835 55275 12841
rect 55217 12832 55229 12835
rect 55088 12804 55229 12832
rect 55088 12792 55094 12804
rect 55217 12801 55229 12804
rect 55263 12801 55275 12835
rect 55217 12795 55275 12801
rect 56410 12792 56416 12844
rect 56468 12832 56474 12844
rect 58345 12835 58403 12841
rect 58345 12832 58357 12835
rect 56468 12804 58357 12832
rect 56468 12792 56474 12804
rect 58345 12801 58357 12804
rect 58391 12801 58403 12835
rect 58345 12795 58403 12801
rect 33091 12736 34560 12764
rect 34977 12767 35035 12773
rect 33091 12733 33103 12736
rect 33045 12727 33103 12733
rect 34977 12733 34989 12767
rect 35023 12764 35035 12767
rect 35894 12764 35900 12776
rect 35023 12736 35900 12764
rect 35023 12733 35035 12736
rect 34977 12727 35035 12733
rect 35894 12724 35900 12736
rect 35952 12724 35958 12776
rect 36078 12764 36084 12776
rect 36039 12736 36084 12764
rect 36078 12724 36084 12736
rect 36136 12724 36142 12776
rect 36170 12724 36176 12776
rect 36228 12773 36234 12776
rect 36228 12767 36251 12773
rect 36239 12733 36251 12767
rect 36538 12764 36544 12776
rect 36228 12727 36251 12733
rect 36280 12736 36544 12764
rect 36228 12724 36234 12727
rect 33502 12696 33508 12708
rect 30607 12668 32352 12696
rect 32416 12668 33508 12696
rect 30607 12665 30619 12668
rect 30561 12659 30619 12665
rect 27948 12600 29592 12628
rect 27948 12588 27954 12600
rect 29638 12588 29644 12640
rect 29696 12628 29702 12640
rect 30837 12631 30895 12637
rect 30837 12628 30849 12631
rect 29696 12600 30849 12628
rect 29696 12588 29702 12600
rect 30837 12597 30849 12600
rect 30883 12597 30895 12631
rect 32324 12628 32352 12668
rect 33502 12656 33508 12668
rect 33560 12656 33566 12708
rect 36280 12696 36308 12736
rect 36538 12724 36544 12736
rect 36596 12764 36602 12776
rect 37458 12764 37464 12776
rect 36596 12736 37464 12764
rect 36596 12724 36602 12736
rect 37458 12724 37464 12736
rect 37516 12724 37522 12776
rect 37573 12767 37631 12773
rect 37573 12764 37585 12767
rect 37568 12733 37585 12764
rect 37619 12733 37631 12767
rect 37568 12727 37631 12733
rect 38013 12767 38071 12773
rect 38013 12733 38025 12767
rect 38059 12764 38071 12767
rect 38838 12764 38844 12776
rect 38059 12736 38844 12764
rect 38059 12733 38071 12736
rect 38013 12727 38071 12733
rect 34992 12668 36308 12696
rect 34992 12628 35020 12668
rect 35158 12628 35164 12640
rect 32324 12600 35020 12628
rect 35119 12600 35164 12628
rect 30837 12591 30895 12597
rect 35158 12588 35164 12600
rect 35216 12588 35222 12640
rect 36170 12588 36176 12640
rect 36228 12628 36234 12640
rect 37568 12628 37596 12727
rect 38838 12724 38844 12736
rect 38896 12724 38902 12776
rect 40589 12767 40647 12773
rect 40589 12733 40601 12767
rect 40635 12733 40647 12767
rect 40589 12727 40647 12733
rect 40604 12696 40632 12727
rect 40678 12724 40684 12776
rect 40736 12764 40742 12776
rect 41969 12767 42027 12773
rect 41969 12764 41981 12767
rect 40736 12736 41981 12764
rect 40736 12724 40742 12736
rect 41969 12733 41981 12736
rect 42015 12733 42027 12767
rect 41969 12727 42027 12733
rect 42061 12767 42119 12773
rect 42061 12733 42073 12767
rect 42107 12733 42119 12767
rect 42061 12727 42119 12733
rect 44177 12767 44235 12773
rect 44177 12733 44189 12767
rect 44223 12733 44235 12767
rect 44358 12764 44364 12776
rect 44319 12736 44364 12764
rect 44177 12727 44235 12733
rect 42076 12696 42104 12727
rect 43438 12696 43444 12708
rect 40604 12668 43444 12696
rect 43438 12656 43444 12668
rect 43496 12656 43502 12708
rect 36228 12600 37596 12628
rect 44192 12628 44220 12727
rect 44358 12724 44364 12736
rect 44416 12724 44422 12776
rect 45370 12764 45376 12776
rect 45331 12736 45376 12764
rect 45370 12724 45376 12736
rect 45428 12724 45434 12776
rect 46753 12767 46811 12773
rect 46753 12733 46765 12767
rect 46799 12733 46811 12767
rect 46753 12727 46811 12733
rect 46768 12696 46796 12727
rect 47026 12724 47032 12776
rect 47084 12764 47090 12776
rect 47121 12767 47179 12773
rect 47121 12764 47133 12767
rect 47084 12736 47133 12764
rect 47084 12724 47090 12736
rect 47121 12733 47133 12736
rect 47167 12733 47179 12767
rect 48130 12764 48136 12776
rect 48091 12736 48136 12764
rect 47121 12727 47179 12733
rect 48130 12724 48136 12736
rect 48188 12724 48194 12776
rect 50246 12764 50252 12776
rect 50207 12736 50252 12764
rect 50246 12724 50252 12736
rect 50304 12724 50310 12776
rect 50341 12767 50399 12773
rect 50341 12733 50353 12767
rect 50387 12764 50399 12767
rect 51074 12764 51080 12776
rect 50387 12736 51080 12764
rect 50387 12733 50399 12736
rect 50341 12727 50399 12733
rect 51074 12724 51080 12736
rect 51132 12724 51138 12776
rect 51626 12724 51632 12776
rect 51684 12764 51690 12776
rect 53285 12767 53343 12773
rect 53285 12764 53297 12767
rect 51684 12736 53297 12764
rect 51684 12724 51690 12736
rect 53285 12733 53297 12736
rect 53331 12733 53343 12767
rect 53285 12727 53343 12733
rect 53653 12767 53711 12773
rect 53653 12733 53665 12767
rect 53699 12733 53711 12767
rect 55306 12764 55312 12776
rect 55267 12736 55312 12764
rect 53653 12727 53711 12733
rect 48038 12696 48044 12708
rect 46768 12668 48044 12696
rect 48038 12656 48044 12668
rect 48096 12656 48102 12708
rect 50062 12696 50068 12708
rect 48240 12668 50068 12696
rect 48240 12628 48268 12668
rect 50062 12656 50068 12668
rect 50120 12696 50126 12708
rect 50890 12696 50896 12708
rect 50120 12668 50896 12696
rect 50120 12656 50126 12668
rect 50890 12656 50896 12668
rect 50948 12656 50954 12708
rect 52730 12656 52736 12708
rect 52788 12696 52794 12708
rect 53668 12696 53696 12727
rect 55306 12724 55312 12736
rect 55364 12724 55370 12776
rect 55677 12767 55735 12773
rect 55677 12733 55689 12767
rect 55723 12733 55735 12767
rect 55677 12727 55735 12733
rect 52788 12668 53696 12696
rect 55692 12696 55720 12727
rect 55766 12724 55772 12776
rect 55824 12764 55830 12776
rect 55824 12736 55869 12764
rect 55824 12724 55830 12736
rect 58434 12724 58440 12776
rect 58492 12764 58498 12776
rect 58621 12767 58679 12773
rect 58621 12764 58633 12767
rect 58492 12736 58633 12764
rect 58492 12724 58498 12736
rect 58621 12733 58633 12736
rect 58667 12733 58679 12767
rect 58621 12727 58679 12733
rect 56134 12696 56140 12708
rect 55692 12668 56140 12696
rect 52788 12656 52794 12668
rect 56134 12656 56140 12668
rect 56192 12656 56198 12708
rect 59722 12628 59728 12640
rect 44192 12600 48268 12628
rect 59683 12600 59728 12628
rect 36228 12588 36234 12600
rect 59722 12588 59728 12600
rect 59780 12588 59786 12640
rect 1104 12538 62192 12560
rect 1104 12486 21344 12538
rect 21396 12486 21408 12538
rect 21460 12486 21472 12538
rect 21524 12486 21536 12538
rect 21588 12486 41707 12538
rect 41759 12486 41771 12538
rect 41823 12486 41835 12538
rect 41887 12486 41899 12538
rect 41951 12486 62192 12538
rect 1104 12464 62192 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 9858 12424 9864 12436
rect 2832 12396 9864 12424
rect 2832 12384 2838 12396
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 9953 12427 10011 12433
rect 9953 12393 9965 12427
rect 9999 12393 10011 12427
rect 9953 12387 10011 12393
rect 5353 12359 5411 12365
rect 5353 12325 5365 12359
rect 5399 12356 5411 12359
rect 5810 12356 5816 12368
rect 5399 12328 5816 12356
rect 5399 12325 5411 12328
rect 5353 12319 5411 12325
rect 5810 12316 5816 12328
rect 5868 12316 5874 12368
rect 6454 12316 6460 12368
rect 6512 12356 6518 12368
rect 7929 12359 7987 12365
rect 6512 12328 7604 12356
rect 6512 12316 6518 12328
rect 5997 12291 6055 12297
rect 5997 12257 6009 12291
rect 6043 12257 6055 12291
rect 6362 12288 6368 12300
rect 6323 12260 6368 12288
rect 5997 12251 6055 12257
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 5905 12223 5963 12229
rect 5905 12220 5917 12223
rect 5684 12192 5917 12220
rect 5684 12180 5690 12192
rect 5905 12189 5917 12192
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 5920 12084 5948 12183
rect 6012 12152 6040 12251
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 6564 12297 6592 12328
rect 6549 12291 6607 12297
rect 6549 12257 6561 12291
rect 6595 12257 6607 12291
rect 7466 12288 7472 12300
rect 7427 12260 7472 12288
rect 6549 12251 6607 12257
rect 7466 12248 7472 12260
rect 7524 12248 7530 12300
rect 6822 12180 6828 12232
rect 6880 12220 6886 12232
rect 7377 12223 7435 12229
rect 7377 12220 7389 12223
rect 6880 12192 7389 12220
rect 6880 12180 6886 12192
rect 7377 12189 7389 12192
rect 7423 12189 7435 12223
rect 7576 12220 7604 12328
rect 7929 12325 7941 12359
rect 7975 12356 7987 12359
rect 9306 12356 9312 12368
rect 7975 12328 9312 12356
rect 7975 12325 7987 12328
rect 7929 12319 7987 12325
rect 9306 12316 9312 12328
rect 9364 12316 9370 12368
rect 9968 12356 9996 12387
rect 11146 12384 11152 12436
rect 11204 12424 11210 12436
rect 11204 12396 12480 12424
rect 11204 12384 11210 12396
rect 11422 12356 11428 12368
rect 9968 12328 11428 12356
rect 11422 12316 11428 12328
rect 11480 12356 11486 12368
rect 12342 12356 12348 12368
rect 11480 12328 12348 12356
rect 11480 12316 11486 12328
rect 9769 12291 9827 12297
rect 9769 12257 9781 12291
rect 9815 12288 9827 12291
rect 10778 12288 10784 12300
rect 9815 12260 10784 12288
rect 9815 12257 9827 12260
rect 9769 12251 9827 12257
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 11514 12288 11520 12300
rect 11475 12260 11520 12288
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 11882 12288 11888 12300
rect 11843 12260 11888 12288
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 11992 12297 12020 12328
rect 12342 12316 12348 12328
rect 12400 12316 12406 12368
rect 11977 12291 12035 12297
rect 11977 12257 11989 12291
rect 12023 12257 12035 12291
rect 12452 12288 12480 12396
rect 18874 12384 18880 12436
rect 18932 12424 18938 12436
rect 18932 12396 21864 12424
rect 18932 12384 18938 12396
rect 16114 12316 16120 12368
rect 16172 12356 16178 12368
rect 17405 12359 17463 12365
rect 17405 12356 17417 12359
rect 16172 12328 17417 12356
rect 16172 12316 16178 12328
rect 17405 12325 17417 12328
rect 17451 12325 17463 12359
rect 17405 12319 17463 12325
rect 18969 12359 19027 12365
rect 18969 12325 18981 12359
rect 19015 12356 19027 12359
rect 19334 12356 19340 12368
rect 19015 12328 19340 12356
rect 19015 12325 19027 12328
rect 18969 12319 19027 12325
rect 19334 12316 19340 12328
rect 19392 12316 19398 12368
rect 19702 12356 19708 12368
rect 19628 12328 19708 12356
rect 12989 12291 13047 12297
rect 12989 12288 13001 12291
rect 12452 12260 13001 12288
rect 11977 12251 12035 12257
rect 12989 12257 13001 12260
rect 13035 12257 13047 12291
rect 12989 12251 13047 12257
rect 15010 12248 15016 12300
rect 15068 12288 15074 12300
rect 16025 12291 16083 12297
rect 16025 12288 16037 12291
rect 15068 12260 16037 12288
rect 15068 12248 15074 12260
rect 16025 12257 16037 12260
rect 16071 12257 16083 12291
rect 16025 12251 16083 12257
rect 16209 12291 16267 12297
rect 16209 12257 16221 12291
rect 16255 12288 16267 12291
rect 16666 12288 16672 12300
rect 16255 12260 16672 12288
rect 16255 12257 16267 12260
rect 16209 12251 16267 12257
rect 16666 12248 16672 12260
rect 16724 12248 16730 12300
rect 17586 12288 17592 12300
rect 17547 12260 17592 12288
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 17770 12248 17776 12300
rect 17828 12288 17834 12300
rect 19628 12288 19656 12328
rect 19702 12316 19708 12328
rect 19760 12356 19766 12368
rect 21634 12356 21640 12368
rect 19760 12328 21640 12356
rect 19760 12316 19766 12328
rect 21634 12316 21640 12328
rect 21692 12316 21698 12368
rect 19794 12288 19800 12300
rect 17828 12260 19656 12288
rect 19755 12260 19800 12288
rect 17828 12248 17834 12260
rect 19794 12248 19800 12260
rect 19852 12248 19858 12300
rect 19981 12291 20039 12297
rect 19981 12257 19993 12291
rect 20027 12288 20039 12291
rect 21726 12288 21732 12300
rect 20027 12260 21588 12288
rect 21687 12260 21732 12288
rect 20027 12257 20039 12260
rect 19981 12251 20039 12257
rect 7926 12220 7932 12232
rect 7576 12192 7932 12220
rect 7377 12183 7435 12189
rect 7926 12180 7932 12192
rect 7984 12180 7990 12232
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12220 10931 12223
rect 10962 12220 10968 12232
rect 10919 12192 10968 12220
rect 10919 12189 10931 12192
rect 10873 12183 10931 12189
rect 10962 12180 10968 12192
rect 11020 12180 11026 12232
rect 11422 12220 11428 12232
rect 11383 12192 11428 12220
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 12894 12220 12900 12232
rect 12855 12192 12900 12220
rect 12894 12180 12900 12192
rect 12952 12180 12958 12232
rect 16577 12223 16635 12229
rect 16577 12189 16589 12223
rect 16623 12189 16635 12223
rect 16577 12183 16635 12189
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12220 18015 12223
rect 19521 12223 19579 12229
rect 19521 12220 19533 12223
rect 18003 12192 19533 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 19521 12189 19533 12192
rect 19567 12189 19579 12223
rect 19521 12183 19579 12189
rect 20901 12223 20959 12229
rect 20901 12189 20913 12223
rect 20947 12220 20959 12223
rect 21082 12220 21088 12232
rect 20947 12192 21088 12220
rect 20947 12189 20959 12192
rect 20901 12183 20959 12189
rect 7098 12152 7104 12164
rect 6012 12124 7104 12152
rect 7098 12112 7104 12124
rect 7156 12112 7162 12164
rect 7558 12152 7564 12164
rect 7208 12124 7564 12152
rect 7208 12084 7236 12124
rect 7558 12112 7564 12124
rect 7616 12112 7622 12164
rect 13078 12112 13084 12164
rect 13136 12152 13142 12164
rect 16390 12152 16396 12164
rect 13136 12124 16396 12152
rect 13136 12112 13142 12124
rect 16390 12112 16396 12124
rect 16448 12112 16454 12164
rect 16592 12152 16620 12183
rect 21082 12180 21088 12192
rect 21140 12180 21146 12232
rect 21453 12223 21511 12229
rect 21453 12189 21465 12223
rect 21499 12189 21511 12223
rect 21560 12220 21588 12260
rect 21726 12248 21732 12260
rect 21784 12248 21790 12300
rect 21836 12288 21864 12396
rect 22278 12384 22284 12436
rect 22336 12424 22342 12436
rect 23017 12427 23075 12433
rect 23017 12424 23029 12427
rect 22336 12396 23029 12424
rect 22336 12384 22342 12396
rect 23017 12393 23029 12396
rect 23063 12393 23075 12427
rect 23842 12424 23848 12436
rect 23017 12387 23075 12393
rect 23124 12396 23848 12424
rect 23124 12356 23152 12396
rect 23842 12384 23848 12396
rect 23900 12424 23906 12436
rect 24305 12427 24363 12433
rect 23900 12396 23980 12424
rect 23900 12384 23906 12396
rect 22848 12328 23152 12356
rect 23952 12356 23980 12396
rect 24305 12393 24317 12427
rect 24351 12424 24363 12427
rect 24394 12424 24400 12436
rect 24351 12396 24400 12424
rect 24351 12393 24363 12396
rect 24305 12387 24363 12393
rect 24394 12384 24400 12396
rect 24452 12384 24458 12436
rect 30006 12424 30012 12436
rect 24504 12396 30012 12424
rect 24504 12356 24532 12396
rect 30006 12384 30012 12396
rect 30064 12384 30070 12436
rect 30653 12427 30711 12433
rect 30653 12393 30665 12427
rect 30699 12424 30711 12427
rect 41414 12424 41420 12436
rect 30699 12396 41420 12424
rect 30699 12393 30711 12396
rect 30653 12387 30711 12393
rect 41414 12384 41420 12396
rect 41472 12384 41478 12436
rect 49973 12427 50031 12433
rect 43364 12396 49924 12424
rect 29638 12356 29644 12368
rect 23952 12328 24532 12356
rect 29380 12328 29644 12356
rect 22741 12291 22799 12297
rect 22741 12288 22753 12291
rect 21836 12260 22753 12288
rect 22741 12257 22753 12260
rect 22787 12257 22799 12291
rect 22741 12251 22799 12257
rect 21913 12223 21971 12229
rect 21913 12220 21925 12223
rect 21560 12192 21925 12220
rect 21453 12183 21511 12189
rect 21913 12189 21925 12192
rect 21959 12220 21971 12223
rect 22848 12220 22876 12328
rect 22925 12291 22983 12297
rect 22925 12257 22937 12291
rect 22971 12257 22983 12291
rect 22925 12251 22983 12257
rect 21959 12192 22876 12220
rect 22940 12220 22968 12251
rect 23566 12248 23572 12300
rect 23624 12288 23630 12300
rect 24118 12288 24124 12300
rect 23624 12260 24124 12288
rect 23624 12248 23630 12260
rect 24118 12248 24124 12260
rect 24176 12248 24182 12300
rect 25222 12248 25228 12300
rect 25280 12248 25286 12300
rect 25317 12291 25375 12297
rect 25317 12257 25329 12291
rect 25363 12288 25375 12291
rect 25406 12288 25412 12300
rect 25363 12260 25412 12288
rect 25363 12257 25375 12260
rect 25317 12251 25375 12257
rect 25406 12248 25412 12260
rect 25464 12248 25470 12300
rect 26605 12291 26663 12297
rect 26605 12257 26617 12291
rect 26651 12288 26663 12291
rect 26697 12291 26755 12297
rect 26697 12288 26709 12291
rect 26651 12260 26709 12288
rect 26651 12257 26663 12260
rect 26605 12251 26663 12257
rect 26697 12257 26709 12260
rect 26743 12257 26755 12291
rect 26697 12251 26755 12257
rect 26881 12291 26939 12297
rect 26881 12257 26893 12291
rect 26927 12257 26939 12291
rect 26881 12251 26939 12257
rect 27249 12291 27307 12297
rect 27249 12257 27261 12291
rect 27295 12288 27307 12291
rect 28537 12291 28595 12297
rect 28537 12288 28549 12291
rect 27295 12260 28549 12288
rect 27295 12257 27307 12260
rect 27249 12251 27307 12257
rect 28537 12257 28549 12260
rect 28583 12257 28595 12291
rect 28718 12288 28724 12300
rect 28679 12260 28724 12288
rect 28537 12251 28595 12257
rect 23474 12220 23480 12232
rect 22940 12192 23480 12220
rect 21959 12189 21971 12192
rect 21913 12183 21971 12189
rect 21468 12152 21496 12183
rect 23474 12180 23480 12192
rect 23532 12220 23538 12232
rect 24302 12220 24308 12232
rect 23532 12192 24308 12220
rect 23532 12180 23538 12192
rect 24302 12180 24308 12192
rect 24360 12180 24366 12232
rect 25240 12220 25268 12248
rect 26896 12220 26924 12251
rect 28718 12248 28724 12260
rect 28776 12248 28782 12300
rect 28810 12248 28816 12300
rect 28868 12288 28874 12300
rect 29380 12297 29408 12328
rect 29638 12316 29644 12328
rect 29696 12316 29702 12368
rect 30098 12316 30104 12368
rect 30156 12356 30162 12368
rect 30156 12328 30604 12356
rect 30156 12316 30162 12328
rect 28905 12291 28963 12297
rect 28905 12288 28917 12291
rect 28868 12260 28917 12288
rect 28868 12248 28874 12260
rect 28905 12257 28917 12260
rect 28951 12257 28963 12291
rect 28905 12251 28963 12257
rect 29365 12291 29423 12297
rect 29365 12257 29377 12291
rect 29411 12257 29423 12291
rect 29365 12251 29423 12257
rect 29549 12291 29607 12297
rect 29549 12257 29561 12291
rect 29595 12288 29607 12291
rect 30190 12288 30196 12300
rect 29595 12260 30196 12288
rect 29595 12257 29607 12260
rect 29549 12251 29607 12257
rect 30190 12248 30196 12260
rect 30248 12248 30254 12300
rect 30576 12297 30604 12328
rect 30742 12316 30748 12368
rect 30800 12356 30806 12368
rect 30800 12328 30845 12356
rect 30800 12316 30806 12328
rect 31018 12316 31024 12368
rect 31076 12356 31082 12368
rect 31113 12359 31171 12365
rect 31113 12356 31125 12359
rect 31076 12328 31125 12356
rect 31076 12316 31082 12328
rect 31113 12325 31125 12328
rect 31159 12325 31171 12359
rect 31113 12319 31171 12325
rect 32125 12359 32183 12365
rect 32125 12325 32137 12359
rect 32171 12356 32183 12359
rect 32398 12356 32404 12368
rect 32171 12328 32404 12356
rect 32171 12325 32183 12328
rect 32125 12319 32183 12325
rect 32398 12316 32404 12328
rect 32456 12316 32462 12368
rect 32950 12356 32956 12368
rect 32692 12328 32956 12356
rect 30561 12291 30619 12297
rect 30561 12257 30573 12291
rect 30607 12288 30619 12291
rect 30607 12260 31156 12288
rect 30607 12257 30619 12260
rect 30561 12251 30619 12257
rect 28074 12220 28080 12232
rect 25240 12192 26924 12220
rect 28035 12192 28080 12220
rect 28074 12180 28080 12192
rect 28132 12180 28138 12232
rect 30377 12223 30435 12229
rect 30377 12220 30389 12223
rect 28184 12192 30389 12220
rect 16592 12124 21496 12152
rect 21542 12112 21548 12164
rect 21600 12152 21606 12164
rect 22002 12152 22008 12164
rect 21600 12124 22008 12152
rect 21600 12112 21606 12124
rect 22002 12112 22008 12124
rect 22060 12152 22066 12164
rect 22060 12124 23704 12152
rect 22060 12112 22066 12124
rect 23676 12096 23704 12124
rect 24946 12112 24952 12164
rect 25004 12152 25010 12164
rect 28184 12152 28212 12192
rect 30377 12189 30389 12192
rect 30423 12220 30435 12223
rect 30466 12220 30472 12232
rect 30423 12192 30472 12220
rect 30423 12189 30435 12192
rect 30377 12183 30435 12189
rect 30466 12180 30472 12192
rect 30524 12180 30530 12232
rect 25004 12124 28212 12152
rect 25004 12112 25010 12124
rect 28258 12112 28264 12164
rect 28316 12152 28322 12164
rect 31018 12152 31024 12164
rect 28316 12124 31024 12152
rect 28316 12112 28322 12124
rect 31018 12112 31024 12124
rect 31076 12112 31082 12164
rect 31128 12152 31156 12260
rect 32214 12248 32220 12300
rect 32272 12288 32278 12300
rect 32692 12288 32720 12328
rect 32950 12316 32956 12328
rect 33008 12316 33014 12368
rect 36630 12356 36636 12368
rect 33336 12328 36308 12356
rect 36591 12328 36636 12356
rect 32272 12260 32720 12288
rect 32272 12248 32278 12260
rect 32766 12248 32772 12300
rect 32824 12288 32830 12300
rect 32968 12288 32996 12316
rect 33336 12297 33364 12328
rect 33103 12291 33161 12297
rect 33103 12288 33115 12291
rect 32824 12260 32869 12288
rect 32968 12260 33115 12288
rect 32824 12248 32830 12260
rect 33103 12257 33115 12260
rect 33149 12257 33161 12291
rect 33103 12251 33161 12257
rect 33321 12291 33379 12297
rect 33321 12257 33333 12291
rect 33367 12257 33379 12291
rect 34330 12288 34336 12300
rect 34291 12260 34336 12288
rect 33321 12251 33379 12257
rect 34330 12248 34336 12260
rect 34388 12248 34394 12300
rect 34425 12291 34483 12297
rect 34425 12257 34437 12291
rect 34471 12257 34483 12291
rect 36170 12288 36176 12300
rect 36131 12260 36176 12288
rect 34425 12251 34483 12257
rect 31202 12180 31208 12232
rect 31260 12220 31266 12232
rect 32582 12220 32588 12232
rect 31260 12192 32588 12220
rect 31260 12180 31266 12192
rect 32582 12180 32588 12192
rect 32640 12180 32646 12232
rect 32861 12223 32919 12229
rect 32861 12189 32873 12223
rect 32907 12220 32919 12223
rect 33778 12220 33784 12232
rect 32907 12192 33784 12220
rect 32907 12189 32919 12192
rect 32861 12183 32919 12189
rect 33778 12180 33784 12192
rect 33836 12180 33842 12232
rect 33962 12180 33968 12232
rect 34020 12220 34026 12232
rect 34440 12220 34468 12251
rect 36170 12248 36176 12260
rect 36228 12248 36234 12300
rect 36280 12288 36308 12328
rect 36630 12316 36636 12328
rect 36688 12316 36694 12368
rect 41138 12316 41144 12368
rect 41196 12356 41202 12368
rect 43364 12356 43392 12396
rect 44542 12356 44548 12368
rect 41196 12328 43392 12356
rect 44503 12328 44548 12356
rect 41196 12316 41202 12328
rect 41233 12291 41291 12297
rect 36280 12260 39620 12288
rect 34020 12192 34468 12220
rect 34020 12180 34026 12192
rect 34974 12180 34980 12232
rect 35032 12220 35038 12232
rect 36081 12223 36139 12229
rect 36081 12220 36093 12223
rect 35032 12192 36093 12220
rect 35032 12180 35038 12192
rect 36081 12189 36093 12192
rect 36127 12189 36139 12223
rect 36081 12183 36139 12189
rect 36446 12180 36452 12232
rect 36504 12220 36510 12232
rect 37826 12220 37832 12232
rect 36504 12192 37832 12220
rect 36504 12180 36510 12192
rect 37826 12180 37832 12192
rect 37884 12220 37890 12232
rect 38746 12220 38752 12232
rect 37884 12192 38752 12220
rect 37884 12180 37890 12192
rect 38746 12180 38752 12192
rect 38804 12180 38810 12232
rect 39022 12220 39028 12232
rect 38983 12192 39028 12220
rect 39022 12180 39028 12192
rect 39080 12180 39086 12232
rect 39592 12220 39620 12260
rect 41233 12257 41245 12291
rect 41279 12288 41291 12291
rect 41414 12288 41420 12300
rect 41279 12260 41420 12288
rect 41279 12257 41291 12260
rect 41233 12251 41291 12257
rect 41414 12248 41420 12260
rect 41472 12248 41478 12300
rect 41506 12248 41512 12300
rect 41564 12288 41570 12300
rect 41693 12291 41751 12297
rect 41693 12288 41705 12291
rect 41564 12260 41705 12288
rect 41564 12248 41570 12260
rect 41693 12257 41705 12260
rect 41739 12257 41751 12291
rect 42058 12288 42064 12300
rect 41971 12260 42064 12288
rect 41693 12251 41751 12257
rect 42058 12248 42064 12260
rect 42116 12288 42122 12300
rect 42242 12288 42248 12300
rect 42116 12260 42248 12288
rect 42116 12248 42122 12260
rect 42242 12248 42248 12260
rect 42300 12248 42306 12300
rect 43364 12297 43392 12328
rect 44542 12316 44548 12328
rect 44600 12316 44606 12368
rect 47118 12356 47124 12368
rect 47079 12328 47124 12356
rect 47118 12316 47124 12328
rect 47176 12316 47182 12368
rect 49896 12356 49924 12396
rect 49973 12393 49985 12427
rect 50019 12424 50031 12427
rect 53190 12424 53196 12436
rect 50019 12396 53196 12424
rect 50019 12393 50031 12396
rect 49973 12387 50031 12393
rect 50522 12356 50528 12368
rect 49896 12328 50528 12356
rect 50522 12316 50528 12328
rect 50580 12356 50586 12368
rect 52457 12359 52515 12365
rect 50580 12328 51028 12356
rect 50580 12316 50586 12328
rect 43349 12291 43407 12297
rect 43349 12257 43361 12291
rect 43395 12257 43407 12291
rect 45186 12288 45192 12300
rect 45147 12260 45192 12288
rect 43349 12251 43407 12257
rect 45186 12248 45192 12260
rect 45244 12248 45250 12300
rect 45554 12288 45560 12300
rect 45515 12260 45560 12288
rect 45554 12248 45560 12260
rect 45612 12248 45618 12300
rect 45741 12291 45799 12297
rect 45741 12257 45753 12291
rect 45787 12288 45799 12291
rect 45830 12288 45836 12300
rect 45787 12260 45836 12288
rect 45787 12257 45799 12260
rect 45741 12251 45799 12257
rect 45830 12248 45836 12260
rect 45888 12248 45894 12300
rect 46661 12291 46719 12297
rect 46661 12257 46673 12291
rect 46707 12257 46719 12291
rect 46661 12251 46719 12257
rect 41966 12220 41972 12232
rect 39592 12192 41972 12220
rect 41966 12180 41972 12192
rect 42024 12180 42030 12232
rect 42150 12220 42156 12232
rect 42111 12192 42156 12220
rect 42150 12180 42156 12192
rect 42208 12180 42214 12232
rect 44726 12180 44732 12232
rect 44784 12220 44790 12232
rect 45097 12223 45155 12229
rect 45097 12220 45109 12223
rect 44784 12192 45109 12220
rect 44784 12180 44790 12192
rect 45097 12189 45109 12192
rect 45143 12189 45155 12223
rect 46566 12220 46572 12232
rect 46527 12192 46572 12220
rect 45097 12183 45155 12189
rect 46566 12180 46572 12192
rect 46624 12180 46630 12232
rect 34149 12155 34207 12161
rect 34149 12152 34161 12155
rect 31128 12124 34161 12152
rect 34149 12121 34161 12124
rect 34195 12121 34207 12155
rect 34149 12115 34207 12121
rect 43438 12112 43444 12164
rect 43496 12152 43502 12164
rect 43533 12155 43591 12161
rect 43533 12152 43545 12155
rect 43496 12124 43545 12152
rect 43496 12112 43502 12124
rect 43533 12121 43545 12124
rect 43579 12152 43591 12155
rect 43806 12152 43812 12164
rect 43579 12124 43812 12152
rect 43579 12121 43591 12124
rect 43533 12115 43591 12121
rect 43806 12112 43812 12124
rect 43864 12152 43870 12164
rect 46198 12152 46204 12164
rect 43864 12124 46204 12152
rect 43864 12112 43870 12124
rect 46198 12112 46204 12124
rect 46256 12152 46262 12164
rect 46676 12152 46704 12251
rect 48222 12248 48228 12300
rect 48280 12288 48286 12300
rect 49789 12291 49847 12297
rect 49789 12288 49801 12291
rect 48280 12260 49801 12288
rect 48280 12248 48286 12260
rect 49789 12257 49801 12260
rect 49835 12257 49847 12291
rect 50890 12288 50896 12300
rect 50851 12260 50896 12288
rect 49789 12251 49847 12257
rect 50890 12248 50896 12260
rect 50948 12248 50954 12300
rect 51000 12297 51028 12328
rect 52457 12325 52469 12359
rect 52503 12356 52515 12359
rect 52546 12356 52552 12368
rect 52503 12328 52552 12356
rect 52503 12325 52515 12328
rect 52457 12319 52515 12325
rect 52546 12316 52552 12328
rect 52604 12316 52610 12368
rect 50985 12291 51043 12297
rect 50985 12257 50997 12291
rect 51031 12257 51043 12291
rect 50985 12251 51043 12257
rect 51445 12223 51503 12229
rect 51445 12189 51457 12223
rect 51491 12189 51503 12223
rect 52932 12220 52960 12396
rect 53190 12384 53196 12396
rect 53248 12424 53254 12436
rect 55030 12424 55036 12436
rect 53248 12396 55036 12424
rect 53248 12384 53254 12396
rect 55030 12384 55036 12396
rect 55088 12384 55094 12436
rect 54570 12356 54576 12368
rect 54531 12328 54576 12356
rect 54570 12316 54576 12328
rect 54628 12316 54634 12368
rect 54680 12328 55812 12356
rect 53101 12291 53159 12297
rect 53101 12257 53113 12291
rect 53147 12257 53159 12291
rect 53466 12288 53472 12300
rect 53427 12260 53472 12288
rect 53101 12251 53159 12257
rect 53009 12223 53067 12229
rect 53009 12220 53021 12223
rect 52932 12192 53021 12220
rect 51445 12183 51503 12189
rect 53009 12189 53021 12192
rect 53055 12189 53067 12223
rect 53116 12220 53144 12251
rect 53466 12248 53472 12260
rect 53524 12248 53530 12300
rect 53558 12248 53564 12300
rect 53616 12288 53622 12300
rect 53653 12291 53711 12297
rect 53653 12288 53665 12291
rect 53616 12260 53665 12288
rect 53616 12248 53622 12260
rect 53653 12257 53665 12260
rect 53699 12288 53711 12291
rect 54680 12288 54708 12328
rect 55784 12300 55812 12328
rect 55858 12316 55864 12368
rect 55916 12356 55922 12368
rect 55916 12328 58572 12356
rect 55916 12316 55922 12328
rect 53699 12260 54708 12288
rect 53699 12257 53711 12260
rect 53653 12251 53711 12257
rect 55030 12248 55036 12300
rect 55088 12288 55094 12300
rect 55217 12291 55275 12297
rect 55217 12288 55229 12291
rect 55088 12260 55229 12288
rect 55088 12248 55094 12260
rect 55217 12257 55229 12260
rect 55263 12257 55275 12291
rect 55217 12251 55275 12257
rect 55585 12291 55643 12297
rect 55585 12257 55597 12291
rect 55631 12257 55643 12291
rect 55766 12288 55772 12300
rect 55727 12260 55772 12288
rect 55585 12251 55643 12257
rect 53742 12220 53748 12232
rect 53116 12192 53748 12220
rect 53009 12183 53067 12189
rect 46256 12124 46704 12152
rect 51460 12152 51488 12183
rect 53742 12180 53748 12192
rect 53800 12180 53806 12232
rect 55125 12223 55183 12229
rect 55125 12189 55137 12223
rect 55171 12189 55183 12223
rect 55125 12183 55183 12189
rect 55140 12152 55168 12183
rect 51460 12124 55168 12152
rect 46256 12112 46262 12124
rect 55214 12112 55220 12164
rect 55272 12152 55278 12164
rect 55600 12152 55628 12251
rect 55766 12248 55772 12260
rect 55824 12248 55830 12300
rect 58158 12288 58164 12300
rect 58119 12260 58164 12288
rect 58158 12248 58164 12260
rect 58216 12248 58222 12300
rect 58544 12297 58572 12328
rect 58345 12291 58403 12297
rect 58345 12257 58357 12291
rect 58391 12257 58403 12291
rect 58345 12251 58403 12257
rect 58529 12291 58587 12297
rect 58529 12257 58541 12291
rect 58575 12288 58587 12291
rect 59722 12288 59728 12300
rect 58575 12260 59728 12288
rect 58575 12257 58587 12260
rect 58529 12251 58587 12257
rect 56042 12180 56048 12232
rect 56100 12220 56106 12232
rect 58360 12220 58388 12251
rect 59722 12248 59728 12260
rect 59780 12248 59786 12300
rect 59078 12220 59084 12232
rect 56100 12192 59084 12220
rect 56100 12180 56106 12192
rect 59078 12180 59084 12192
rect 59136 12180 59142 12232
rect 55272 12124 55628 12152
rect 57977 12155 58035 12161
rect 55272 12112 55278 12124
rect 57977 12121 57989 12155
rect 58023 12152 58035 12155
rect 58434 12152 58440 12164
rect 58023 12124 58440 12152
rect 58023 12121 58035 12124
rect 57977 12115 58035 12121
rect 58434 12112 58440 12124
rect 58492 12112 58498 12164
rect 5920 12056 7236 12084
rect 7282 12044 7288 12096
rect 7340 12084 7346 12096
rect 8202 12084 8208 12096
rect 7340 12056 8208 12084
rect 7340 12044 7346 12056
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 12986 12044 12992 12096
rect 13044 12084 13050 12096
rect 13173 12087 13231 12093
rect 13173 12084 13185 12087
rect 13044 12056 13185 12084
rect 13044 12044 13050 12056
rect 13173 12053 13185 12056
rect 13219 12053 13231 12087
rect 13173 12047 13231 12053
rect 13354 12044 13360 12096
rect 13412 12084 13418 12096
rect 13538 12084 13544 12096
rect 13412 12056 13544 12084
rect 13412 12044 13418 12056
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 15102 12084 15108 12096
rect 14056 12056 15108 12084
rect 14056 12044 14062 12056
rect 15102 12044 15108 12056
rect 15160 12044 15166 12096
rect 15378 12044 15384 12096
rect 15436 12084 15442 12096
rect 23566 12084 23572 12096
rect 15436 12056 23572 12084
rect 15436 12044 15442 12056
rect 23566 12044 23572 12056
rect 23624 12044 23630 12096
rect 23658 12044 23664 12096
rect 23716 12084 23722 12096
rect 25498 12084 25504 12096
rect 23716 12056 25504 12084
rect 23716 12044 23722 12056
rect 25498 12044 25504 12056
rect 25556 12044 25562 12096
rect 26605 12087 26663 12093
rect 26605 12053 26617 12087
rect 26651 12084 26663 12087
rect 34238 12084 34244 12096
rect 26651 12056 34244 12084
rect 26651 12053 26663 12056
rect 26605 12047 26663 12053
rect 34238 12044 34244 12056
rect 34296 12044 34302 12096
rect 34422 12044 34428 12096
rect 34480 12084 34486 12096
rect 34609 12087 34667 12093
rect 34609 12084 34621 12087
rect 34480 12056 34621 12084
rect 34480 12044 34486 12056
rect 34609 12053 34621 12056
rect 34655 12053 34667 12087
rect 34609 12047 34667 12053
rect 35894 12044 35900 12096
rect 35952 12084 35958 12096
rect 36722 12084 36728 12096
rect 35952 12056 36728 12084
rect 35952 12044 35958 12056
rect 36722 12044 36728 12056
rect 36780 12044 36786 12096
rect 37182 12044 37188 12096
rect 37240 12084 37246 12096
rect 39666 12084 39672 12096
rect 37240 12056 39672 12084
rect 37240 12044 37246 12056
rect 39666 12044 39672 12056
rect 39724 12044 39730 12096
rect 40126 12084 40132 12096
rect 40087 12056 40132 12084
rect 40126 12044 40132 12056
rect 40184 12084 40190 12096
rect 40678 12084 40684 12096
rect 40184 12056 40684 12084
rect 40184 12044 40190 12056
rect 40678 12044 40684 12056
rect 40736 12044 40742 12096
rect 50246 12044 50252 12096
rect 50304 12084 50310 12096
rect 56226 12084 56232 12096
rect 50304 12056 56232 12084
rect 50304 12044 50310 12056
rect 56226 12044 56232 12056
rect 56284 12044 56290 12096
rect 1104 11994 62192 12016
rect 1104 11942 11163 11994
rect 11215 11942 11227 11994
rect 11279 11942 11291 11994
rect 11343 11942 11355 11994
rect 11407 11942 31526 11994
rect 31578 11942 31590 11994
rect 31642 11942 31654 11994
rect 31706 11942 31718 11994
rect 31770 11942 51888 11994
rect 51940 11942 51952 11994
rect 52004 11942 52016 11994
rect 52068 11942 52080 11994
rect 52132 11942 62192 11994
rect 1104 11920 62192 11942
rect 6917 11883 6975 11889
rect 6917 11849 6929 11883
rect 6963 11880 6975 11883
rect 7190 11880 7196 11892
rect 6963 11852 7196 11880
rect 6963 11849 6975 11852
rect 6917 11843 6975 11849
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 13170 11880 13176 11892
rect 7300 11852 13176 11880
rect 7300 11812 7328 11852
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 13262 11840 13268 11892
rect 13320 11880 13326 11892
rect 19886 11880 19892 11892
rect 13320 11852 19892 11880
rect 13320 11840 13326 11852
rect 19886 11840 19892 11852
rect 19944 11840 19950 11892
rect 20070 11880 20076 11892
rect 20031 11852 20076 11880
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 21542 11880 21548 11892
rect 20548 11852 21548 11880
rect 12342 11812 12348 11824
rect 4448 11784 7328 11812
rect 7760 11784 12348 11812
rect 3050 11744 3056 11756
rect 3011 11716 3056 11744
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 3142 11676 3148 11688
rect 3103 11648 3148 11676
rect 3142 11636 3148 11648
rect 3200 11636 3206 11688
rect 4448 11685 4476 11784
rect 4816 11716 7512 11744
rect 4433 11679 4491 11685
rect 4433 11645 4445 11679
rect 4479 11645 4491 11679
rect 4433 11639 4491 11645
rect 3605 11611 3663 11617
rect 3605 11577 3617 11611
rect 3651 11608 3663 11611
rect 4816 11608 4844 11716
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11645 4951 11679
rect 5074 11676 5080 11688
rect 5035 11648 5080 11676
rect 4893 11639 4951 11645
rect 3651 11580 4844 11608
rect 3651 11577 3663 11580
rect 3605 11571 3663 11577
rect 4908 11540 4936 11639
rect 5074 11636 5080 11648
rect 5132 11636 5138 11688
rect 5353 11679 5411 11685
rect 5353 11645 5365 11679
rect 5399 11645 5411 11679
rect 5353 11639 5411 11645
rect 5368 11608 5396 11639
rect 5442 11636 5448 11688
rect 5500 11676 5506 11688
rect 5537 11679 5595 11685
rect 5537 11676 5549 11679
rect 5500 11648 5549 11676
rect 5500 11636 5506 11648
rect 5537 11645 5549 11648
rect 5583 11645 5595 11679
rect 5537 11639 5595 11645
rect 5905 11679 5963 11685
rect 5905 11645 5917 11679
rect 5951 11676 5963 11679
rect 6914 11676 6920 11688
rect 5951 11648 6920 11676
rect 5951 11645 5963 11648
rect 5905 11639 5963 11645
rect 6914 11636 6920 11648
rect 6972 11636 6978 11688
rect 7484 11685 7512 11716
rect 7558 11704 7564 11756
rect 7616 11744 7622 11756
rect 7616 11716 7661 11744
rect 7616 11704 7622 11716
rect 7469 11679 7527 11685
rect 7469 11645 7481 11679
rect 7515 11645 7527 11679
rect 7469 11639 7527 11645
rect 7760 11608 7788 11784
rect 12342 11772 12348 11784
rect 12400 11772 12406 11824
rect 12529 11815 12587 11821
rect 12529 11781 12541 11815
rect 12575 11812 12587 11815
rect 12710 11812 12716 11824
rect 12575 11784 12716 11812
rect 12575 11781 12587 11784
rect 12529 11775 12587 11781
rect 12710 11772 12716 11784
rect 12768 11772 12774 11824
rect 14366 11772 14372 11824
rect 14424 11812 14430 11824
rect 20548 11812 20576 11852
rect 21542 11840 21548 11852
rect 21600 11840 21606 11892
rect 22094 11840 22100 11892
rect 22152 11880 22158 11892
rect 22281 11883 22339 11889
rect 22281 11880 22293 11883
rect 22152 11852 22293 11880
rect 22152 11840 22158 11852
rect 22281 11849 22293 11852
rect 22327 11849 22339 11883
rect 22281 11843 22339 11849
rect 25498 11840 25504 11892
rect 25556 11880 25562 11892
rect 25556 11852 32168 11880
rect 25556 11840 25562 11852
rect 23385 11815 23443 11821
rect 23385 11812 23397 11815
rect 14424 11784 20576 11812
rect 20640 11784 23397 11812
rect 14424 11772 14430 11784
rect 7926 11744 7932 11756
rect 7839 11716 7932 11744
rect 7926 11704 7932 11716
rect 7984 11744 7990 11756
rect 11238 11744 11244 11756
rect 7984 11716 11244 11744
rect 7984 11704 7990 11716
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 11514 11744 11520 11756
rect 11475 11716 11520 11744
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 12434 11704 12440 11756
rect 12492 11744 12498 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12492 11716 13001 11744
rect 12492 11704 12498 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 13354 11704 13360 11756
rect 13412 11744 13418 11756
rect 13541 11747 13599 11753
rect 13541 11744 13553 11747
rect 13412 11716 13553 11744
rect 13412 11704 13418 11716
rect 13541 11713 13553 11716
rect 13587 11744 13599 11747
rect 13630 11744 13636 11756
rect 13587 11716 13636 11744
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 15010 11744 15016 11756
rect 14292 11716 15016 11744
rect 7837 11679 7895 11685
rect 7837 11645 7849 11679
rect 7883 11676 7895 11679
rect 8018 11676 8024 11688
rect 7883 11648 8024 11676
rect 7883 11645 7895 11648
rect 7837 11639 7895 11645
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 8202 11636 8208 11688
rect 8260 11676 8266 11688
rect 8849 11679 8907 11685
rect 8849 11676 8861 11679
rect 8260 11648 8861 11676
rect 8260 11636 8266 11648
rect 8849 11645 8861 11648
rect 8895 11645 8907 11679
rect 9030 11676 9036 11688
rect 8943 11648 9036 11676
rect 8849 11639 8907 11645
rect 9030 11636 9036 11648
rect 9088 11676 9094 11688
rect 10965 11679 11023 11685
rect 9088 11648 9812 11676
rect 9088 11636 9094 11648
rect 5368 11580 7788 11608
rect 9125 11543 9183 11549
rect 9125 11540 9137 11543
rect 4908 11512 9137 11540
rect 9125 11509 9137 11512
rect 9171 11509 9183 11543
rect 9784 11540 9812 11648
rect 10965 11645 10977 11679
rect 11011 11645 11023 11679
rect 10965 11639 11023 11645
rect 10980 11608 11008 11639
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11112 11648 11157 11676
rect 11112 11636 11118 11648
rect 11330 11636 11336 11688
rect 11388 11676 11394 11688
rect 13081 11679 13139 11685
rect 13081 11676 13093 11679
rect 11388 11648 13093 11676
rect 11388 11636 11394 11648
rect 13081 11645 13093 11648
rect 13127 11645 13139 11679
rect 13081 11639 13139 11645
rect 13262 11636 13268 11688
rect 13320 11676 13326 11688
rect 13449 11679 13507 11685
rect 13449 11676 13461 11679
rect 13320 11648 13461 11676
rect 13320 11636 13326 11648
rect 13449 11645 13461 11648
rect 13495 11645 13507 11679
rect 13449 11639 13507 11645
rect 14292 11608 14320 11716
rect 15010 11704 15016 11716
rect 15068 11744 15074 11756
rect 15068 11716 15332 11744
rect 15068 11704 15074 11716
rect 14918 11676 14924 11688
rect 14879 11648 14924 11676
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 15304 11685 15332 11716
rect 15378 11704 15384 11756
rect 15436 11744 15442 11756
rect 18417 11747 18475 11753
rect 15436 11716 15481 11744
rect 15436 11704 15442 11716
rect 18417 11713 18429 11747
rect 18463 11744 18475 11747
rect 20254 11744 20260 11756
rect 18463 11716 20260 11744
rect 18463 11713 18475 11716
rect 18417 11707 18475 11713
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 15289 11679 15347 11685
rect 15289 11645 15301 11679
rect 15335 11645 15347 11679
rect 15289 11639 15347 11645
rect 16206 11636 16212 11688
rect 16264 11676 16270 11688
rect 16485 11679 16543 11685
rect 16485 11676 16497 11679
rect 16264 11648 16497 11676
rect 16264 11636 16270 11648
rect 16485 11645 16497 11648
rect 16531 11645 16543 11679
rect 16485 11639 16543 11645
rect 16761 11679 16819 11685
rect 16761 11645 16773 11679
rect 16807 11645 16819 11679
rect 16761 11639 16819 11645
rect 17129 11679 17187 11685
rect 17129 11645 17141 11679
rect 17175 11676 17187 11679
rect 18693 11679 18751 11685
rect 18693 11676 18705 11679
rect 17175 11648 18705 11676
rect 17175 11645 17187 11648
rect 17129 11639 17187 11645
rect 18693 11645 18705 11648
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 14458 11608 14464 11620
rect 10980 11580 14320 11608
rect 14419 11580 14464 11608
rect 14458 11568 14464 11580
rect 14516 11568 14522 11620
rect 14550 11568 14556 11620
rect 14608 11608 14614 11620
rect 16577 11611 16635 11617
rect 16577 11608 16589 11611
rect 14608 11580 16589 11608
rect 14608 11568 14614 11580
rect 16577 11577 16589 11580
rect 16623 11577 16635 11611
rect 16776 11608 16804 11639
rect 19702 11636 19708 11688
rect 19760 11676 19766 11688
rect 20640 11685 20668 11784
rect 23385 11781 23397 11784
rect 23431 11781 23443 11815
rect 23385 11775 23443 11781
rect 23750 11772 23756 11824
rect 23808 11812 23814 11824
rect 23845 11815 23903 11821
rect 23845 11812 23857 11815
rect 23808 11784 23857 11812
rect 23808 11772 23814 11784
rect 23845 11781 23857 11784
rect 23891 11812 23903 11815
rect 28350 11812 28356 11824
rect 23891 11784 28356 11812
rect 23891 11781 23903 11784
rect 23845 11775 23903 11781
rect 28350 11772 28356 11784
rect 28408 11772 28414 11824
rect 30190 11772 30196 11824
rect 30248 11812 30254 11824
rect 30248 11784 31616 11812
rect 30248 11772 30254 11784
rect 20806 11704 20812 11756
rect 20864 11744 20870 11756
rect 21082 11744 21088 11756
rect 20864 11716 20944 11744
rect 21043 11716 21088 11744
rect 20864 11704 20870 11716
rect 20625 11679 20683 11685
rect 20625 11676 20637 11679
rect 19760 11648 20637 11676
rect 19760 11636 19766 11648
rect 20625 11645 20637 11648
rect 20671 11645 20683 11679
rect 20625 11639 20683 11645
rect 20717 11679 20775 11685
rect 20717 11645 20729 11679
rect 20763 11676 20775 11679
rect 20916 11676 20944 11716
rect 21082 11704 21088 11716
rect 21140 11704 21146 11756
rect 21726 11704 21732 11756
rect 21784 11744 21790 11756
rect 26881 11747 26939 11753
rect 21784 11716 23704 11744
rect 21784 11704 21790 11716
rect 20993 11679 21051 11685
rect 20993 11676 21005 11679
rect 20763 11648 20852 11676
rect 20916 11648 21005 11676
rect 20763 11645 20775 11648
rect 20717 11639 20775 11645
rect 17494 11608 17500 11620
rect 16776 11580 17500 11608
rect 16577 11571 16635 11577
rect 17494 11568 17500 11580
rect 17552 11568 17558 11620
rect 18782 11608 18788 11620
rect 18743 11580 18788 11608
rect 18782 11568 18788 11580
rect 18840 11568 18846 11620
rect 19153 11611 19211 11617
rect 19153 11577 19165 11611
rect 19199 11608 19211 11611
rect 19334 11608 19340 11620
rect 19199 11580 19340 11608
rect 19199 11577 19211 11580
rect 19153 11571 19211 11577
rect 19334 11568 19340 11580
rect 19392 11568 19398 11620
rect 12802 11540 12808 11552
rect 9784 11512 12808 11540
rect 9125 11503 9183 11509
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 15746 11500 15752 11552
rect 15804 11540 15810 11552
rect 16298 11540 16304 11552
rect 15804 11512 16304 11540
rect 15804 11500 15810 11512
rect 16298 11500 16304 11512
rect 16356 11500 16362 11552
rect 18601 11543 18659 11549
rect 18601 11509 18613 11543
rect 18647 11540 18659 11543
rect 20622 11540 20628 11552
rect 18647 11512 20628 11540
rect 18647 11509 18659 11512
rect 18601 11503 18659 11509
rect 20622 11500 20628 11512
rect 20680 11500 20686 11552
rect 20824 11540 20852 11648
rect 20993 11645 21005 11648
rect 21039 11645 21051 11679
rect 20993 11639 21051 11645
rect 22189 11679 22247 11685
rect 22189 11645 22201 11679
rect 22235 11676 22247 11679
rect 23474 11676 23480 11688
rect 22235 11648 23480 11676
rect 22235 11645 22247 11648
rect 22189 11639 22247 11645
rect 23474 11636 23480 11648
rect 23532 11636 23538 11688
rect 23676 11685 23704 11716
rect 26881 11713 26893 11747
rect 26927 11744 26939 11747
rect 27338 11744 27344 11756
rect 26927 11716 27344 11744
rect 26927 11713 26939 11716
rect 26881 11707 26939 11713
rect 27338 11704 27344 11716
rect 27396 11704 27402 11756
rect 27614 11744 27620 11756
rect 27448 11716 27620 11744
rect 23661 11679 23719 11685
rect 23661 11645 23673 11679
rect 23707 11676 23719 11679
rect 24026 11676 24032 11688
rect 23707 11648 24032 11676
rect 23707 11645 23719 11648
rect 23661 11639 23719 11645
rect 24026 11636 24032 11648
rect 24084 11636 24090 11688
rect 24762 11676 24768 11688
rect 24723 11648 24768 11676
rect 24762 11636 24768 11648
rect 24820 11636 24826 11688
rect 25774 11636 25780 11688
rect 25832 11676 25838 11688
rect 25869 11679 25927 11685
rect 25869 11676 25881 11679
rect 25832 11648 25881 11676
rect 25832 11636 25838 11648
rect 25869 11645 25881 11648
rect 25915 11645 25927 11679
rect 25869 11639 25927 11645
rect 26142 11636 26148 11688
rect 26200 11676 26206 11688
rect 26786 11676 26792 11688
rect 26200 11648 26792 11676
rect 26200 11636 26206 11648
rect 26786 11636 26792 11648
rect 26844 11636 26850 11688
rect 27448 11685 27476 11716
rect 27614 11704 27620 11716
rect 27672 11704 27678 11756
rect 27890 11744 27896 11756
rect 27724 11716 27896 11744
rect 27724 11685 27752 11716
rect 27890 11704 27896 11716
rect 27948 11704 27954 11756
rect 28074 11744 28080 11756
rect 28035 11716 28080 11744
rect 28074 11704 28080 11716
rect 28132 11704 28138 11756
rect 28368 11744 28396 11772
rect 30561 11747 30619 11753
rect 28368 11716 30512 11744
rect 27433 11679 27491 11685
rect 27433 11645 27445 11679
rect 27479 11645 27491 11679
rect 27433 11639 27491 11645
rect 27525 11679 27583 11685
rect 27525 11645 27537 11679
rect 27571 11645 27583 11679
rect 27525 11639 27583 11645
rect 27709 11679 27767 11685
rect 27709 11645 27721 11679
rect 27755 11645 27767 11679
rect 27709 11639 27767 11645
rect 20898 11568 20904 11620
rect 20956 11608 20962 11620
rect 22005 11611 22063 11617
rect 22005 11608 22017 11611
rect 20956 11580 22017 11608
rect 20956 11568 20962 11580
rect 22005 11577 22017 11580
rect 22051 11577 22063 11611
rect 22005 11571 22063 11577
rect 23385 11611 23443 11617
rect 23385 11577 23397 11611
rect 23431 11608 23443 11611
rect 27338 11608 27344 11620
rect 23431 11580 27344 11608
rect 23431 11577 23443 11580
rect 23385 11571 23443 11577
rect 22462 11540 22468 11552
rect 20824 11512 22468 11540
rect 22462 11500 22468 11512
rect 22520 11500 22526 11552
rect 24964 11549 24992 11580
rect 27338 11568 27344 11580
rect 27396 11568 27402 11620
rect 27540 11608 27568 11639
rect 27798 11636 27804 11688
rect 27856 11676 27862 11688
rect 28261 11679 28319 11685
rect 28261 11676 28273 11679
rect 27856 11648 28273 11676
rect 27856 11636 27862 11648
rect 28261 11645 28273 11648
rect 28307 11676 28319 11679
rect 30190 11676 30196 11688
rect 28307 11648 29960 11676
rect 30151 11648 30196 11676
rect 28307 11645 28319 11648
rect 28261 11639 28319 11645
rect 29822 11608 29828 11620
rect 27540 11580 29828 11608
rect 29822 11568 29828 11580
rect 29880 11568 29886 11620
rect 24949 11543 25007 11549
rect 24949 11509 24961 11543
rect 24995 11509 25007 11543
rect 24949 11503 25007 11509
rect 25314 11500 25320 11552
rect 25372 11540 25378 11552
rect 25961 11543 26019 11549
rect 25961 11540 25973 11543
rect 25372 11512 25973 11540
rect 25372 11500 25378 11512
rect 25961 11509 25973 11512
rect 26007 11509 26019 11543
rect 25961 11503 26019 11509
rect 26050 11500 26056 11552
rect 26108 11540 26114 11552
rect 27982 11540 27988 11552
rect 26108 11512 27988 11540
rect 26108 11500 26114 11512
rect 27982 11500 27988 11512
rect 28040 11500 28046 11552
rect 29932 11540 29960 11648
rect 30190 11636 30196 11648
rect 30248 11636 30254 11688
rect 30484 11676 30512 11716
rect 30561 11713 30573 11747
rect 30607 11744 30619 11747
rect 30742 11744 30748 11756
rect 30607 11716 30748 11744
rect 30607 11713 30619 11716
rect 30561 11707 30619 11713
rect 30742 11704 30748 11716
rect 30800 11704 30806 11756
rect 31588 11753 31616 11784
rect 32140 11753 32168 11852
rect 32398 11840 32404 11892
rect 32456 11880 32462 11892
rect 32456 11852 34284 11880
rect 32456 11840 32462 11852
rect 34256 11812 34284 11852
rect 34330 11840 34336 11892
rect 34388 11880 34394 11892
rect 35161 11883 35219 11889
rect 35161 11880 35173 11883
rect 34388 11852 35173 11880
rect 34388 11840 34394 11852
rect 35161 11849 35173 11852
rect 35207 11849 35219 11883
rect 38930 11880 38936 11892
rect 35161 11843 35219 11849
rect 36372 11852 38936 11880
rect 36372 11812 36400 11852
rect 38930 11840 38936 11852
rect 38988 11880 38994 11892
rect 40126 11880 40132 11892
rect 38988 11852 40132 11880
rect 38988 11840 38994 11852
rect 40126 11840 40132 11852
rect 40184 11840 40190 11892
rect 45186 11840 45192 11892
rect 45244 11880 45250 11892
rect 46385 11883 46443 11889
rect 46385 11880 46397 11883
rect 45244 11852 46397 11880
rect 45244 11840 45250 11852
rect 46385 11849 46397 11852
rect 46431 11849 46443 11883
rect 46385 11843 46443 11849
rect 49694 11840 49700 11892
rect 49752 11880 49758 11892
rect 49752 11852 52684 11880
rect 49752 11840 49758 11852
rect 33152 11784 34192 11812
rect 34256 11784 36400 11812
rect 31573 11747 31631 11753
rect 31573 11713 31585 11747
rect 31619 11713 31631 11747
rect 31573 11707 31631 11713
rect 32125 11747 32183 11753
rect 32125 11713 32137 11747
rect 32171 11744 32183 11747
rect 32171 11716 32536 11744
rect 32171 11713 32183 11716
rect 32125 11707 32183 11713
rect 32214 11676 32220 11688
rect 30484 11648 32220 11676
rect 32214 11636 32220 11648
rect 32272 11636 32278 11688
rect 32398 11676 32404 11688
rect 32359 11648 32404 11676
rect 32398 11636 32404 11648
rect 32456 11636 32462 11688
rect 32508 11676 32536 11716
rect 32582 11704 32588 11756
rect 32640 11744 32646 11756
rect 33152 11744 33180 11784
rect 33686 11744 33692 11756
rect 32640 11716 33180 11744
rect 33244 11716 33692 11744
rect 32640 11704 32646 11716
rect 33244 11676 33272 11716
rect 33686 11704 33692 11716
rect 33744 11704 33750 11756
rect 33962 11744 33968 11756
rect 33923 11716 33968 11744
rect 33962 11704 33968 11716
rect 34020 11704 34026 11756
rect 34164 11744 34192 11784
rect 37366 11772 37372 11824
rect 37424 11812 37430 11824
rect 41598 11812 41604 11824
rect 37424 11784 41604 11812
rect 37424 11772 37430 11784
rect 41598 11772 41604 11784
rect 41656 11772 41662 11824
rect 43714 11772 43720 11824
rect 43772 11812 43778 11824
rect 43772 11784 45232 11812
rect 43772 11772 43778 11784
rect 34164 11716 34744 11744
rect 32508 11648 33272 11676
rect 33502 11636 33508 11688
rect 33560 11676 33566 11688
rect 33597 11679 33655 11685
rect 33597 11676 33609 11679
rect 33560 11648 33609 11676
rect 33560 11636 33566 11648
rect 33597 11645 33609 11648
rect 33643 11676 33655 11679
rect 34146 11676 34152 11688
rect 33643 11648 34152 11676
rect 33643 11645 33655 11648
rect 33597 11639 33655 11645
rect 34146 11636 34152 11648
rect 34204 11636 34210 11688
rect 34716 11676 34744 11716
rect 34790 11704 34796 11756
rect 34848 11744 34854 11756
rect 41230 11744 41236 11756
rect 34848 11716 41236 11744
rect 34848 11704 34854 11716
rect 41230 11704 41236 11716
rect 41288 11704 41294 11756
rect 41414 11704 41420 11756
rect 41472 11744 41478 11756
rect 41877 11747 41935 11753
rect 41877 11744 41889 11747
rect 41472 11716 41889 11744
rect 41472 11704 41478 11716
rect 41877 11713 41889 11716
rect 41923 11713 41935 11747
rect 41877 11707 41935 11713
rect 41966 11704 41972 11756
rect 42024 11744 42030 11756
rect 44085 11747 44143 11753
rect 44085 11744 44097 11747
rect 42024 11716 44097 11744
rect 42024 11704 42030 11716
rect 44085 11713 44097 11716
rect 44131 11713 44143 11747
rect 44085 11707 44143 11713
rect 44358 11704 44364 11756
rect 44416 11744 44422 11756
rect 45097 11747 45155 11753
rect 45097 11744 45109 11747
rect 44416 11716 45109 11744
rect 44416 11704 44422 11716
rect 45097 11713 45109 11716
rect 45143 11713 45155 11747
rect 45204 11744 45232 11784
rect 45278 11772 45284 11824
rect 45336 11812 45342 11824
rect 46658 11812 46664 11824
rect 45336 11784 46664 11812
rect 45336 11772 45342 11784
rect 46658 11772 46664 11784
rect 46716 11772 46722 11824
rect 48593 11815 48651 11821
rect 48593 11781 48605 11815
rect 48639 11812 48651 11815
rect 49234 11812 49240 11824
rect 48639 11784 49240 11812
rect 48639 11781 48651 11784
rect 48593 11775 48651 11781
rect 49234 11772 49240 11784
rect 49292 11772 49298 11824
rect 51994 11812 52000 11824
rect 51955 11784 52000 11812
rect 51994 11772 52000 11784
rect 52052 11772 52058 11824
rect 52656 11812 52684 11852
rect 52914 11840 52920 11892
rect 52972 11880 52978 11892
rect 55858 11880 55864 11892
rect 52972 11852 55864 11880
rect 52972 11840 52978 11852
rect 55858 11840 55864 11852
rect 55916 11840 55922 11892
rect 60458 11880 60464 11892
rect 56704 11852 60464 11880
rect 56042 11812 56048 11824
rect 52656 11784 56048 11812
rect 46109 11747 46167 11753
rect 46109 11744 46121 11747
rect 45204 11716 46121 11744
rect 45097 11707 45155 11713
rect 46109 11713 46121 11716
rect 46155 11713 46167 11747
rect 46109 11707 46167 11713
rect 46290 11704 46296 11756
rect 46348 11744 46354 11756
rect 52656 11753 52684 11784
rect 56042 11772 56048 11784
rect 56100 11772 56106 11824
rect 52641 11747 52699 11753
rect 46348 11716 52592 11744
rect 46348 11704 46354 11716
rect 35069 11679 35127 11685
rect 35069 11676 35081 11679
rect 34716 11648 35081 11676
rect 35069 11645 35081 11648
rect 35115 11676 35127 11679
rect 35710 11676 35716 11688
rect 35115 11648 35716 11676
rect 35115 11645 35127 11648
rect 35069 11639 35127 11645
rect 35710 11636 35716 11648
rect 35768 11636 35774 11688
rect 36357 11679 36415 11685
rect 36357 11645 36369 11679
rect 36403 11676 36415 11679
rect 36446 11676 36452 11688
rect 36403 11648 36452 11676
rect 36403 11645 36415 11648
rect 36357 11639 36415 11645
rect 36446 11636 36452 11648
rect 36504 11636 36510 11688
rect 36630 11676 36636 11688
rect 36591 11648 36636 11676
rect 36630 11636 36636 11648
rect 36688 11636 36694 11688
rect 36722 11636 36728 11688
rect 36780 11676 36786 11688
rect 37090 11676 37096 11688
rect 36780 11648 37096 11676
rect 36780 11636 36786 11648
rect 37090 11636 37096 11648
rect 37148 11676 37154 11688
rect 41138 11676 41144 11688
rect 37148 11648 41144 11676
rect 37148 11636 37154 11648
rect 41138 11636 41144 11648
rect 41196 11636 41202 11688
rect 41601 11679 41659 11685
rect 41601 11645 41613 11679
rect 41647 11676 41659 11679
rect 42334 11676 42340 11688
rect 41647 11648 42340 11676
rect 41647 11645 41659 11648
rect 41601 11639 41659 11645
rect 42334 11636 42340 11648
rect 42392 11676 42398 11688
rect 42392 11648 42564 11676
rect 42392 11636 42398 11648
rect 30009 11611 30067 11617
rect 30009 11577 30021 11611
rect 30055 11608 30067 11611
rect 30650 11608 30656 11620
rect 30055 11580 30656 11608
rect 30055 11577 30067 11580
rect 30009 11571 30067 11577
rect 30650 11568 30656 11580
rect 30708 11568 30714 11620
rect 32766 11608 32772 11620
rect 30760 11580 32772 11608
rect 30760 11540 30788 11580
rect 32766 11568 32772 11580
rect 32824 11568 32830 11620
rect 33413 11611 33471 11617
rect 33413 11577 33425 11611
rect 33459 11608 33471 11611
rect 34790 11608 34796 11620
rect 33459 11580 34796 11608
rect 33459 11577 33471 11580
rect 33413 11571 33471 11577
rect 34790 11568 34796 11580
rect 34848 11568 34854 11620
rect 34885 11611 34943 11617
rect 34885 11577 34897 11611
rect 34931 11577 34943 11611
rect 41414 11608 41420 11620
rect 34885 11571 34943 11577
rect 37568 11580 41420 11608
rect 29932 11512 30788 11540
rect 30834 11500 30840 11552
rect 30892 11540 30898 11552
rect 33962 11540 33968 11552
rect 30892 11512 33968 11540
rect 30892 11500 30898 11512
rect 33962 11500 33968 11512
rect 34020 11500 34026 11552
rect 34900 11540 34928 11571
rect 37568 11540 37596 11580
rect 41414 11568 41420 11580
rect 41472 11568 41478 11620
rect 42536 11608 42564 11648
rect 42610 11636 42616 11688
rect 42668 11676 42674 11688
rect 44637 11679 44695 11685
rect 44637 11676 44649 11679
rect 42668 11648 44649 11676
rect 42668 11636 42674 11648
rect 44637 11645 44649 11648
rect 44683 11645 44695 11679
rect 44637 11639 44695 11645
rect 44913 11679 44971 11685
rect 44913 11645 44925 11679
rect 44959 11645 44971 11679
rect 46198 11676 46204 11688
rect 46159 11648 46204 11676
rect 44913 11639 44971 11645
rect 42886 11608 42892 11620
rect 42536 11580 42892 11608
rect 42886 11568 42892 11580
rect 42944 11568 42950 11620
rect 34900 11512 37596 11540
rect 37642 11500 37648 11552
rect 37700 11540 37706 11552
rect 37737 11543 37795 11549
rect 37737 11540 37749 11543
rect 37700 11512 37749 11540
rect 37700 11500 37706 11512
rect 37737 11509 37749 11512
rect 37783 11509 37795 11543
rect 37737 11503 37795 11509
rect 42242 11500 42248 11552
rect 42300 11540 42306 11552
rect 43162 11540 43168 11552
rect 42300 11512 43168 11540
rect 42300 11500 42306 11512
rect 43162 11500 43168 11512
rect 43220 11500 43226 11552
rect 44928 11540 44956 11639
rect 46198 11636 46204 11648
rect 46256 11636 46262 11688
rect 48774 11676 48780 11688
rect 48735 11648 48780 11676
rect 48774 11636 48780 11648
rect 48832 11636 48838 11688
rect 49145 11679 49203 11685
rect 49145 11645 49157 11679
rect 49191 11645 49203 11679
rect 49145 11639 49203 11645
rect 49237 11679 49295 11685
rect 49237 11645 49249 11679
rect 49283 11676 49295 11679
rect 49694 11676 49700 11688
rect 49283 11648 49700 11676
rect 49283 11645 49295 11648
rect 49237 11639 49295 11645
rect 45186 11568 45192 11620
rect 45244 11608 45250 11620
rect 48682 11608 48688 11620
rect 45244 11580 48688 11608
rect 45244 11568 45250 11580
rect 48682 11568 48688 11580
rect 48740 11568 48746 11620
rect 49160 11608 49188 11639
rect 49694 11636 49700 11648
rect 49752 11636 49758 11688
rect 50522 11676 50528 11688
rect 50483 11648 50528 11676
rect 50522 11636 50528 11648
rect 50580 11636 50586 11688
rect 51626 11636 51632 11688
rect 51684 11676 51690 11688
rect 52564 11685 52592 11716
rect 52641 11713 52653 11747
rect 52687 11713 52699 11747
rect 52641 11707 52699 11713
rect 54297 11747 54355 11753
rect 54297 11713 54309 11747
rect 54343 11744 54355 11747
rect 55306 11744 55312 11756
rect 54343 11716 55312 11744
rect 54343 11713 54355 11716
rect 54297 11707 54355 11713
rect 55306 11704 55312 11716
rect 55364 11704 55370 11756
rect 56704 11744 56732 11852
rect 60458 11840 60464 11852
rect 60516 11840 60522 11892
rect 55876 11716 56732 11744
rect 52181 11679 52239 11685
rect 52181 11676 52193 11679
rect 51684 11648 52193 11676
rect 51684 11636 51690 11648
rect 52181 11645 52193 11648
rect 52227 11645 52239 11679
rect 52181 11639 52239 11645
rect 52549 11679 52607 11685
rect 52549 11645 52561 11679
rect 52595 11676 52607 11679
rect 53190 11676 53196 11688
rect 52595 11648 53196 11676
rect 52595 11645 52607 11648
rect 52549 11639 52607 11645
rect 53190 11636 53196 11648
rect 53248 11676 53254 11688
rect 55876 11685 55904 11716
rect 56778 11704 56784 11756
rect 56836 11744 56842 11756
rect 57977 11747 58035 11753
rect 57977 11744 57989 11747
rect 56836 11716 57989 11744
rect 56836 11704 56842 11716
rect 57977 11713 57989 11716
rect 58023 11713 58035 11747
rect 57977 11707 58035 11713
rect 53745 11679 53803 11685
rect 53745 11676 53757 11679
rect 53248 11648 53757 11676
rect 53248 11636 53254 11648
rect 53745 11645 53757 11648
rect 53791 11645 53803 11679
rect 53745 11639 53803 11645
rect 53837 11679 53895 11685
rect 53837 11645 53849 11679
rect 53883 11645 53895 11679
rect 53837 11639 53895 11645
rect 55861 11679 55919 11685
rect 55861 11645 55873 11679
rect 55907 11645 55919 11679
rect 56226 11676 56232 11688
rect 56187 11648 56232 11676
rect 55861 11639 55919 11645
rect 50614 11608 50620 11620
rect 49160 11580 50620 11608
rect 49160 11540 49188 11580
rect 50614 11568 50620 11580
rect 50672 11568 50678 11620
rect 44928 11512 49188 11540
rect 49970 11500 49976 11552
rect 50028 11540 50034 11552
rect 50522 11540 50528 11552
rect 50028 11512 50528 11540
rect 50028 11500 50034 11512
rect 50522 11500 50528 11512
rect 50580 11500 50586 11552
rect 50709 11543 50767 11549
rect 50709 11509 50721 11543
rect 50755 11540 50767 11543
rect 51074 11540 51080 11552
rect 50755 11512 51080 11540
rect 50755 11509 50767 11512
rect 50709 11503 50767 11509
rect 51074 11500 51080 11512
rect 51132 11540 51138 11552
rect 52362 11540 52368 11552
rect 51132 11512 52368 11540
rect 51132 11500 51138 11512
rect 52362 11500 52368 11512
rect 52420 11540 52426 11552
rect 53852 11540 53880 11639
rect 56226 11636 56232 11648
rect 56284 11636 56290 11688
rect 56321 11679 56379 11685
rect 56321 11645 56333 11679
rect 56367 11676 56379 11679
rect 56594 11676 56600 11688
rect 56367 11648 56600 11676
rect 56367 11645 56379 11648
rect 56321 11639 56379 11645
rect 56594 11636 56600 11648
rect 56652 11636 56658 11688
rect 57330 11636 57336 11688
rect 57388 11676 57394 11688
rect 57701 11679 57759 11685
rect 57701 11676 57713 11679
rect 57388 11648 57713 11676
rect 57388 11636 57394 11648
rect 57701 11645 57713 11648
rect 57747 11645 57759 11679
rect 57701 11639 57759 11645
rect 55401 11611 55459 11617
rect 55401 11577 55413 11611
rect 55447 11608 55459 11611
rect 56686 11608 56692 11620
rect 55447 11580 56692 11608
rect 55447 11577 55459 11580
rect 55401 11571 55459 11577
rect 56686 11568 56692 11580
rect 56744 11568 56750 11620
rect 54662 11540 54668 11552
rect 52420 11512 54668 11540
rect 52420 11500 52426 11512
rect 54662 11500 54668 11512
rect 54720 11500 54726 11552
rect 56226 11500 56232 11552
rect 56284 11540 56290 11552
rect 59081 11543 59139 11549
rect 59081 11540 59093 11543
rect 56284 11512 59093 11540
rect 56284 11500 56290 11512
rect 59081 11509 59093 11512
rect 59127 11509 59139 11543
rect 59081 11503 59139 11509
rect 1104 11450 62192 11472
rect 1104 11398 21344 11450
rect 21396 11398 21408 11450
rect 21460 11398 21472 11450
rect 21524 11398 21536 11450
rect 21588 11398 41707 11450
rect 41759 11398 41771 11450
rect 41823 11398 41835 11450
rect 41887 11398 41899 11450
rect 41951 11398 62192 11450
rect 1104 11376 62192 11398
rect 5074 11336 5080 11348
rect 3160 11308 5080 11336
rect 3160 11277 3188 11308
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 7484 11308 13124 11336
rect 3145 11271 3203 11277
rect 3145 11237 3157 11271
rect 3191 11237 3203 11271
rect 6914 11268 6920 11280
rect 6875 11240 6920 11268
rect 3145 11231 3203 11237
rect 6914 11228 6920 11240
rect 6972 11228 6978 11280
rect 2593 11203 2651 11209
rect 2593 11169 2605 11203
rect 2639 11169 2651 11203
rect 2593 11163 2651 11169
rect 2608 11132 2636 11163
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 2832 11172 2877 11200
rect 2832 11160 2838 11172
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 7484 11209 7512 11308
rect 11330 11268 11336 11280
rect 9692 11240 11100 11268
rect 11291 11240 11336 11268
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4028 11172 4445 11200
rect 4028 11160 4034 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 7469 11203 7527 11209
rect 7469 11169 7481 11203
rect 7515 11169 7527 11203
rect 7469 11163 7527 11169
rect 7745 11203 7803 11209
rect 7745 11169 7757 11203
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 7929 11203 7987 11209
rect 7929 11169 7941 11203
rect 7975 11200 7987 11203
rect 9030 11200 9036 11212
rect 7975 11172 9036 11200
rect 7975 11169 7987 11172
rect 7929 11163 7987 11169
rect 3050 11132 3056 11144
rect 2608 11104 3056 11132
rect 3050 11092 3056 11104
rect 3108 11132 3114 11144
rect 4706 11132 4712 11144
rect 3108 11104 4476 11132
rect 4667 11104 4712 11132
rect 3108 11092 3114 11104
rect 4448 11076 4476 11104
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 6822 11132 6828 11144
rect 5828 11104 6828 11132
rect 4430 11024 4436 11076
rect 4488 11024 4494 11076
rect 5534 11024 5540 11076
rect 5592 11064 5598 11076
rect 5828 11073 5856 11104
rect 6822 11092 6828 11104
rect 6880 11132 6886 11144
rect 7760 11132 7788 11163
rect 9030 11160 9036 11172
rect 9088 11160 9094 11212
rect 9692 11209 9720 11240
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11169 9735 11203
rect 10778 11200 10784 11212
rect 10739 11172 10784 11200
rect 9677 11163 9735 11169
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 10873 11203 10931 11209
rect 10873 11169 10885 11203
rect 10919 11200 10931 11203
rect 10962 11200 10968 11212
rect 10919 11172 10968 11200
rect 10919 11169 10931 11172
rect 10873 11163 10931 11169
rect 6880 11104 7788 11132
rect 6880 11092 6886 11104
rect 5813 11067 5871 11073
rect 5813 11064 5825 11067
rect 5592 11036 5825 11064
rect 5592 11024 5598 11036
rect 5813 11033 5825 11036
rect 5859 11033 5871 11067
rect 5813 11027 5871 11033
rect 7466 11024 7472 11076
rect 7524 11064 7530 11076
rect 9861 11067 9919 11073
rect 9861 11064 9873 11067
rect 7524 11036 9873 11064
rect 7524 11024 7530 11036
rect 9861 11033 9873 11036
rect 9907 11064 9919 11067
rect 10888 11064 10916 11163
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 11072 11200 11100 11240
rect 11330 11228 11336 11240
rect 11388 11228 11394 11280
rect 13096 11268 13124 11308
rect 13170 11296 13176 11348
rect 13228 11336 13234 11348
rect 21082 11336 21088 11348
rect 13228 11308 17356 11336
rect 13228 11296 13234 11308
rect 14366 11268 14372 11280
rect 13096 11240 14372 11268
rect 14366 11228 14372 11240
rect 14424 11228 14430 11280
rect 14918 11228 14924 11280
rect 14976 11268 14982 11280
rect 17328 11277 17356 11308
rect 17420 11308 21088 11336
rect 15841 11271 15899 11277
rect 15841 11268 15853 11271
rect 14976 11240 15853 11268
rect 14976 11228 14982 11240
rect 15841 11237 15853 11240
rect 15887 11237 15899 11271
rect 15841 11231 15899 11237
rect 17313 11271 17371 11277
rect 17313 11237 17325 11271
rect 17359 11237 17371 11271
rect 17313 11231 17371 11237
rect 13998 11200 14004 11212
rect 11072 11172 14004 11200
rect 13998 11160 14004 11172
rect 14056 11160 14062 11212
rect 14090 11160 14096 11212
rect 14148 11200 14154 11212
rect 15289 11203 15347 11209
rect 15289 11200 15301 11203
rect 14148 11172 15301 11200
rect 14148 11160 14154 11172
rect 15289 11169 15301 11172
rect 15335 11169 15347 11203
rect 15289 11163 15347 11169
rect 15381 11203 15439 11209
rect 15381 11169 15393 11203
rect 15427 11200 15439 11203
rect 16022 11200 16028 11212
rect 15427 11172 16028 11200
rect 15427 11169 15439 11172
rect 15381 11163 15439 11169
rect 16022 11160 16028 11172
rect 16080 11160 16086 11212
rect 12158 11092 12164 11144
rect 12216 11132 12222 11144
rect 12437 11135 12495 11141
rect 12216 11104 12261 11132
rect 12216 11092 12222 11104
rect 12437 11101 12449 11135
rect 12483 11132 12495 11135
rect 15102 11132 15108 11144
rect 12483 11104 15108 11132
rect 12483 11101 12495 11104
rect 12437 11095 12495 11101
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 15194 11092 15200 11144
rect 15252 11132 15258 11144
rect 17420 11132 17448 11308
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 21634 11296 21640 11348
rect 21692 11336 21698 11348
rect 24397 11339 24455 11345
rect 24397 11336 24409 11339
rect 21692 11308 24409 11336
rect 21692 11296 21698 11308
rect 24397 11305 24409 11308
rect 24443 11336 24455 11339
rect 28445 11339 28503 11345
rect 28445 11336 28457 11339
rect 24443 11308 25360 11336
rect 24443 11305 24455 11308
rect 24397 11299 24455 11305
rect 18230 11228 18236 11280
rect 18288 11268 18294 11280
rect 18693 11271 18751 11277
rect 18693 11268 18705 11271
rect 18288 11240 18705 11268
rect 18288 11228 18294 11240
rect 18693 11237 18705 11240
rect 18739 11237 18751 11271
rect 18693 11231 18751 11237
rect 18782 11228 18788 11280
rect 18840 11268 18846 11280
rect 18840 11240 19840 11268
rect 18840 11228 18846 11240
rect 17497 11203 17555 11209
rect 17497 11169 17509 11203
rect 17543 11169 17555 11203
rect 19334 11200 19340 11212
rect 19295 11172 19340 11200
rect 17497 11163 17555 11169
rect 15252 11104 17448 11132
rect 15252 11092 15258 11104
rect 9907 11036 10916 11064
rect 9907 11033 9919 11036
rect 9861 11027 9919 11033
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 13725 11067 13783 11073
rect 13725 11064 13737 11067
rect 13504 11036 13737 11064
rect 13504 11024 13510 11036
rect 13725 11033 13737 11036
rect 13771 11064 13783 11067
rect 16114 11064 16120 11076
rect 13771 11036 16120 11064
rect 13771 11033 13783 11036
rect 13725 11027 13783 11033
rect 16114 11024 16120 11036
rect 16172 11024 16178 11076
rect 17512 11008 17540 11163
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 19702 11200 19708 11212
rect 19663 11172 19708 11200
rect 19702 11160 19708 11172
rect 19760 11160 19766 11212
rect 19812 11209 19840 11240
rect 20622 11228 20628 11280
rect 20680 11268 20686 11280
rect 21453 11271 21511 11277
rect 21453 11268 21465 11271
rect 20680 11240 21465 11268
rect 20680 11228 20686 11240
rect 21453 11237 21465 11240
rect 21499 11237 21511 11271
rect 21453 11231 21511 11237
rect 19797 11203 19855 11209
rect 19797 11169 19809 11203
rect 19843 11169 19855 11203
rect 19797 11163 19855 11169
rect 19886 11160 19892 11212
rect 19944 11200 19950 11212
rect 20993 11203 21051 11209
rect 20993 11200 21005 11203
rect 19944 11172 21005 11200
rect 19944 11160 19950 11172
rect 20993 11169 21005 11172
rect 21039 11200 21051 11203
rect 21468 11200 21496 11231
rect 22557 11203 22615 11209
rect 21039 11172 21404 11200
rect 21468 11172 21680 11200
rect 21039 11169 21051 11172
rect 20993 11163 21051 11169
rect 17865 11135 17923 11141
rect 17865 11101 17877 11135
rect 17911 11132 17923 11135
rect 19242 11132 19248 11144
rect 17911 11104 19248 11132
rect 17911 11101 17923 11104
rect 17865 11095 17923 11101
rect 19242 11092 19248 11104
rect 19300 11092 19306 11144
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11132 19487 11135
rect 19610 11132 19616 11144
rect 19475 11104 19616 11132
rect 19475 11101 19487 11104
rect 19429 11095 19487 11101
rect 19610 11092 19616 11104
rect 19668 11092 19674 11144
rect 20254 11092 20260 11144
rect 20312 11132 20318 11144
rect 20898 11132 20904 11144
rect 20312 11104 20904 11132
rect 20312 11092 20318 11104
rect 20898 11092 20904 11104
rect 20956 11092 20962 11144
rect 21376 11064 21404 11172
rect 21652 11132 21680 11172
rect 22557 11169 22569 11203
rect 22603 11200 22615 11203
rect 22646 11200 22652 11212
rect 22603 11172 22652 11200
rect 22603 11169 22615 11172
rect 22557 11163 22615 11169
rect 22646 11160 22652 11172
rect 22704 11160 22710 11212
rect 23109 11203 23167 11209
rect 23109 11169 23121 11203
rect 23155 11169 23167 11203
rect 23290 11200 23296 11212
rect 23251 11172 23296 11200
rect 23109 11163 23167 11169
rect 23124 11132 23152 11163
rect 23290 11160 23296 11172
rect 23348 11160 23354 11212
rect 24210 11200 24216 11212
rect 24171 11172 24216 11200
rect 24210 11160 24216 11172
rect 24268 11160 24274 11212
rect 25332 11209 25360 11308
rect 26804 11308 28457 11336
rect 26804 11277 26832 11308
rect 28445 11305 28457 11308
rect 28491 11305 28503 11339
rect 29822 11336 29828 11348
rect 29783 11308 29828 11336
rect 28445 11299 28503 11305
rect 29822 11296 29828 11308
rect 29880 11296 29886 11348
rect 30926 11296 30932 11348
rect 30984 11336 30990 11348
rect 31110 11336 31116 11348
rect 30984 11308 31116 11336
rect 30984 11296 30990 11308
rect 31110 11296 31116 11308
rect 31168 11296 31174 11348
rect 32306 11336 32312 11348
rect 32219 11308 32312 11336
rect 32306 11296 32312 11308
rect 32364 11336 32370 11348
rect 32364 11308 40172 11336
rect 32364 11296 32370 11308
rect 26789 11271 26847 11277
rect 26789 11237 26801 11271
rect 26835 11237 26847 11271
rect 26789 11231 26847 11237
rect 27154 11228 27160 11280
rect 27212 11268 27218 11280
rect 28169 11271 28227 11277
rect 28169 11268 28181 11271
rect 27212 11240 28181 11268
rect 27212 11228 27218 11240
rect 28169 11237 28181 11240
rect 28215 11237 28227 11271
rect 28169 11231 28227 11237
rect 28258 11228 28264 11280
rect 28316 11268 28322 11280
rect 29549 11271 29607 11277
rect 28316 11240 28488 11268
rect 28316 11228 28322 11240
rect 25317 11203 25375 11209
rect 25317 11169 25329 11203
rect 25363 11200 25375 11203
rect 26050 11200 26056 11212
rect 25363 11172 26056 11200
rect 25363 11169 25375 11172
rect 25317 11163 25375 11169
rect 26050 11160 26056 11172
rect 26108 11160 26114 11212
rect 26881 11203 26939 11209
rect 26881 11169 26893 11203
rect 26927 11200 26939 11203
rect 27614 11200 27620 11212
rect 26927 11172 27620 11200
rect 26927 11169 26939 11172
rect 26881 11163 26939 11169
rect 27614 11160 27620 11172
rect 27672 11160 27678 11212
rect 27890 11200 27896 11212
rect 27724 11172 27896 11200
rect 27724 11132 27752 11172
rect 27890 11160 27896 11172
rect 27948 11160 27954 11212
rect 28350 11200 28356 11212
rect 28311 11172 28356 11200
rect 28350 11160 28356 11172
rect 28408 11160 28414 11212
rect 21652 11104 27752 11132
rect 27798 11092 27804 11144
rect 27856 11132 27862 11144
rect 28460 11132 28488 11240
rect 29549 11237 29561 11271
rect 29595 11268 29607 11271
rect 29595 11240 33364 11268
rect 29595 11237 29607 11240
rect 29549 11231 29607 11237
rect 28994 11160 29000 11212
rect 29052 11200 29058 11212
rect 29733 11203 29791 11209
rect 29733 11200 29745 11203
rect 29052 11172 29745 11200
rect 29052 11160 29058 11172
rect 29733 11169 29745 11172
rect 29779 11200 29791 11203
rect 30190 11200 30196 11212
rect 29779 11172 30196 11200
rect 29779 11169 29791 11172
rect 29733 11163 29791 11169
rect 30190 11160 30196 11172
rect 30248 11160 30254 11212
rect 30466 11160 30472 11212
rect 30524 11200 30530 11212
rect 30929 11203 30987 11209
rect 30929 11200 30941 11203
rect 30524 11172 30941 11200
rect 30524 11160 30530 11172
rect 30929 11169 30941 11172
rect 30975 11169 30987 11203
rect 30929 11163 30987 11169
rect 32125 11203 32183 11209
rect 32125 11169 32137 11203
rect 32171 11169 32183 11203
rect 33336 11200 33364 11240
rect 34238 11228 34244 11280
rect 34296 11268 34302 11280
rect 40144 11268 40172 11308
rect 40494 11296 40500 11348
rect 40552 11336 40558 11348
rect 40589 11339 40647 11345
rect 40589 11336 40601 11339
rect 40552 11308 40601 11336
rect 40552 11296 40558 11308
rect 40589 11305 40601 11308
rect 40635 11305 40647 11339
rect 40589 11299 40647 11305
rect 41414 11296 41420 11348
rect 41472 11336 41478 11348
rect 47486 11336 47492 11348
rect 41472 11308 47492 11336
rect 41472 11296 41478 11308
rect 47486 11296 47492 11308
rect 47544 11336 47550 11348
rect 47544 11308 49924 11336
rect 47544 11296 47550 11308
rect 34296 11240 37872 11268
rect 40144 11240 44036 11268
rect 34296 11228 34302 11240
rect 33336 11172 33916 11200
rect 32125 11163 32183 11169
rect 32140 11132 32168 11163
rect 27856 11104 32168 11132
rect 33229 11135 33287 11141
rect 27856 11092 27862 11104
rect 33229 11101 33241 11135
rect 33275 11101 33287 11135
rect 33502 11132 33508 11144
rect 33463 11104 33508 11132
rect 33229 11095 33287 11101
rect 21726 11064 21732 11076
rect 21376 11036 21732 11064
rect 21726 11024 21732 11036
rect 21784 11024 21790 11076
rect 25501 11067 25559 11073
rect 25501 11033 25513 11067
rect 25547 11064 25559 11067
rect 28994 11064 29000 11076
rect 25547 11036 29000 11064
rect 25547 11033 25559 11036
rect 25501 11027 25559 11033
rect 28994 11024 29000 11036
rect 29052 11024 29058 11076
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 10870 10996 10876 11008
rect 9732 10968 10876 10996
rect 9732 10956 9738 10968
rect 10870 10956 10876 10968
rect 10928 10996 10934 11008
rect 12434 10996 12440 11008
rect 10928 10968 12440 10996
rect 10928 10956 10934 10968
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 17494 10996 17500 11008
rect 17407 10968 17500 10996
rect 17494 10956 17500 10968
rect 17552 10996 17558 11008
rect 22554 10996 22560 11008
rect 17552 10968 22560 10996
rect 17552 10956 17558 10968
rect 22554 10956 22560 10968
rect 22612 10956 22618 11008
rect 23382 10956 23388 11008
rect 23440 10996 23446 11008
rect 26605 10999 26663 11005
rect 23440 10968 23485 10996
rect 23440 10956 23446 10968
rect 26605 10965 26617 10999
rect 26651 10996 26663 10999
rect 26694 10996 26700 11008
rect 26651 10968 26700 10996
rect 26651 10965 26663 10968
rect 26605 10959 26663 10965
rect 26694 10956 26700 10968
rect 26752 10956 26758 11008
rect 27062 10996 27068 11008
rect 27023 10968 27068 10996
rect 27062 10956 27068 10968
rect 27120 10956 27126 11008
rect 33244 10996 33272 11095
rect 33502 11092 33508 11104
rect 33560 11092 33566 11144
rect 33888 11132 33916 11172
rect 33962 11160 33968 11212
rect 34020 11200 34026 11212
rect 34885 11203 34943 11209
rect 34885 11200 34897 11203
rect 34020 11172 34897 11200
rect 34020 11160 34026 11172
rect 34885 11169 34897 11172
rect 34931 11200 34943 11203
rect 35066 11200 35072 11212
rect 34931 11172 35072 11200
rect 34931 11169 34943 11172
rect 34885 11163 34943 11169
rect 35066 11160 35072 11172
rect 35124 11160 35130 11212
rect 36262 11200 36268 11212
rect 36223 11172 36268 11200
rect 36262 11160 36268 11172
rect 36320 11160 36326 11212
rect 36538 11160 36544 11212
rect 36596 11200 36602 11212
rect 36633 11203 36691 11209
rect 36633 11200 36645 11203
rect 36596 11172 36645 11200
rect 36596 11160 36602 11172
rect 36633 11169 36645 11172
rect 36679 11169 36691 11203
rect 36633 11163 36691 11169
rect 36814 11160 36820 11212
rect 36872 11200 36878 11212
rect 37743 11203 37801 11209
rect 37743 11200 37755 11203
rect 36872 11172 37755 11200
rect 36872 11160 36878 11172
rect 37743 11169 37755 11172
rect 37789 11169 37801 11203
rect 37844 11200 37872 11240
rect 41414 11200 41420 11212
rect 37844 11172 41420 11200
rect 37743 11163 37801 11169
rect 41414 11160 41420 11172
rect 41472 11160 41478 11212
rect 41785 11203 41843 11209
rect 41785 11169 41797 11203
rect 41831 11200 41843 11203
rect 41877 11203 41935 11209
rect 41877 11200 41889 11203
rect 41831 11172 41889 11200
rect 41831 11169 41843 11172
rect 41785 11163 41843 11169
rect 41877 11169 41889 11172
rect 41923 11169 41935 11203
rect 41877 11163 41935 11169
rect 42061 11203 42119 11209
rect 42061 11169 42073 11203
rect 42107 11169 42119 11203
rect 42061 11163 42119 11169
rect 42429 11203 42487 11209
rect 42429 11169 42441 11203
rect 42475 11200 42487 11203
rect 42610 11200 42616 11212
rect 42475 11172 42616 11200
rect 42475 11169 42487 11172
rect 42429 11163 42487 11169
rect 34974 11132 34980 11144
rect 33888 11104 34980 11132
rect 34974 11092 34980 11104
rect 35032 11092 35038 11144
rect 36725 11135 36783 11141
rect 36725 11101 36737 11135
rect 36771 11132 36783 11135
rect 36771 11104 37688 11132
rect 36771 11101 36783 11104
rect 36725 11095 36783 11101
rect 36081 11067 36139 11073
rect 36081 11033 36093 11067
rect 36127 11064 36139 11067
rect 36630 11064 36636 11076
rect 36127 11036 36636 11064
rect 36127 11033 36139 11036
rect 36081 11027 36139 11033
rect 36630 11024 36636 11036
rect 36688 11024 36694 11076
rect 33594 10996 33600 11008
rect 33244 10968 33600 10996
rect 33594 10956 33600 10968
rect 33652 10996 33658 11008
rect 34882 10996 34888 11008
rect 33652 10968 34888 10996
rect 33652 10956 33658 10968
rect 34882 10956 34888 10968
rect 34940 10996 34946 11008
rect 36446 10996 36452 11008
rect 34940 10968 36452 10996
rect 34940 10956 34946 10968
rect 36446 10956 36452 10968
rect 36504 10956 36510 11008
rect 37660 10996 37688 11104
rect 38746 11092 38752 11144
rect 38804 11132 38810 11144
rect 39206 11132 39212 11144
rect 38804 11104 39212 11132
rect 38804 11092 38810 11104
rect 39206 11092 39212 11104
rect 39264 11092 39270 11144
rect 39482 11132 39488 11144
rect 39443 11104 39488 11132
rect 39482 11092 39488 11104
rect 39540 11092 39546 11144
rect 41322 11092 41328 11144
rect 41380 11132 41386 11144
rect 42076 11132 42104 11163
rect 42610 11160 42616 11172
rect 42668 11160 42674 11212
rect 43162 11160 43168 11212
rect 43220 11200 43226 11212
rect 43625 11203 43683 11209
rect 43625 11200 43637 11203
rect 43220 11172 43637 11200
rect 43220 11160 43226 11172
rect 43625 11169 43637 11172
rect 43671 11169 43683 11203
rect 43625 11163 43683 11169
rect 43717 11203 43775 11209
rect 43717 11169 43729 11203
rect 43763 11200 43775 11203
rect 43806 11200 43812 11212
rect 43763 11172 43812 11200
rect 43763 11169 43775 11172
rect 43717 11163 43775 11169
rect 43806 11160 43812 11172
rect 43864 11160 43870 11212
rect 44008 11200 44036 11240
rect 44082 11228 44088 11280
rect 44140 11268 44146 11280
rect 44177 11271 44235 11277
rect 44177 11268 44189 11271
rect 44140 11240 44189 11268
rect 44140 11228 44146 11240
rect 44177 11237 44189 11240
rect 44223 11237 44235 11271
rect 48038 11268 48044 11280
rect 47999 11240 48044 11268
rect 44177 11231 44235 11237
rect 48038 11228 48044 11240
rect 48096 11228 48102 11280
rect 47581 11203 47639 11209
rect 47581 11200 47593 11203
rect 44008 11172 47593 11200
rect 47581 11169 47593 11172
rect 47627 11169 47639 11203
rect 47581 11163 47639 11169
rect 48961 11203 49019 11209
rect 48961 11169 48973 11203
rect 49007 11200 49019 11203
rect 49050 11200 49056 11212
rect 49007 11172 49056 11200
rect 49007 11169 49019 11172
rect 48961 11163 49019 11169
rect 49050 11160 49056 11172
rect 49108 11160 49114 11212
rect 49234 11200 49240 11212
rect 49195 11172 49240 11200
rect 49234 11160 49240 11172
rect 49292 11160 49298 11212
rect 49896 11200 49924 11308
rect 51534 11296 51540 11348
rect 51592 11336 51598 11348
rect 53101 11339 53159 11345
rect 51592 11308 53052 11336
rect 51592 11296 51598 11308
rect 50614 11268 50620 11280
rect 50575 11240 50620 11268
rect 50614 11228 50620 11240
rect 50672 11228 50678 11280
rect 53024 11268 53052 11308
rect 53101 11305 53113 11339
rect 53147 11336 53159 11339
rect 53190 11336 53196 11348
rect 53147 11308 53196 11336
rect 53147 11305 53159 11308
rect 53101 11299 53159 11305
rect 53190 11296 53196 11308
rect 53248 11296 53254 11348
rect 53300 11308 55260 11336
rect 53300 11268 53328 11308
rect 53024 11240 53328 11268
rect 53742 11228 53748 11280
rect 53800 11268 53806 11280
rect 55125 11271 55183 11277
rect 55125 11268 55137 11271
rect 53800 11240 55137 11268
rect 53800 11228 53806 11240
rect 55125 11237 55137 11240
rect 55171 11237 55183 11271
rect 55125 11231 55183 11237
rect 51994 11200 52000 11212
rect 49896 11172 51856 11200
rect 51955 11172 52000 11200
rect 44818 11132 44824 11144
rect 41380 11104 44824 11132
rect 41380 11092 41386 11104
rect 44818 11092 44824 11104
rect 44876 11092 44882 11144
rect 45005 11135 45063 11141
rect 45005 11101 45017 11135
rect 45051 11132 45063 11135
rect 45186 11132 45192 11144
rect 45051 11104 45192 11132
rect 45051 11101 45063 11104
rect 45005 11095 45063 11101
rect 45186 11092 45192 11104
rect 45244 11092 45250 11144
rect 45281 11135 45339 11141
rect 45281 11101 45293 11135
rect 45327 11132 45339 11135
rect 46106 11132 46112 11144
rect 45327 11104 46112 11132
rect 45327 11101 45339 11104
rect 45281 11095 45339 11101
rect 46106 11092 46112 11104
rect 46164 11092 46170 11144
rect 47486 11132 47492 11144
rect 47447 11104 47492 11132
rect 47486 11092 47492 11104
rect 47544 11092 47550 11144
rect 51534 11092 51540 11144
rect 51592 11132 51598 11144
rect 51721 11135 51779 11141
rect 51721 11132 51733 11135
rect 51592 11104 51733 11132
rect 51592 11092 51598 11104
rect 51721 11101 51733 11104
rect 51767 11101 51779 11135
rect 51828 11132 51856 11172
rect 51994 11160 52000 11172
rect 52052 11160 52058 11212
rect 54662 11200 54668 11212
rect 54623 11172 54668 11200
rect 54662 11160 54668 11172
rect 54720 11160 54726 11212
rect 55232 11200 55260 11308
rect 56318 11296 56324 11348
rect 56376 11336 56382 11348
rect 57977 11339 58035 11345
rect 57977 11336 57989 11339
rect 56376 11308 57989 11336
rect 56376 11296 56382 11308
rect 57977 11305 57989 11308
rect 58023 11305 58035 11339
rect 59078 11336 59084 11348
rect 59039 11308 59084 11336
rect 57977 11299 58035 11305
rect 59078 11296 59084 11308
rect 59136 11296 59142 11348
rect 56413 11203 56471 11209
rect 56413 11200 56425 11203
rect 55232 11172 56425 11200
rect 56413 11169 56425 11172
rect 56459 11169 56471 11203
rect 56686 11200 56692 11212
rect 56647 11172 56692 11200
rect 56413 11163 56471 11169
rect 51828 11104 54524 11132
rect 51721 11095 51779 11101
rect 37921 11067 37979 11073
rect 37921 11064 37933 11067
rect 37844 11036 37933 11064
rect 37844 10996 37872 11036
rect 37921 11033 37933 11036
rect 37967 11064 37979 11067
rect 38838 11064 38844 11076
rect 37967 11036 38844 11064
rect 37967 11033 37979 11036
rect 37921 11027 37979 11033
rect 38838 11024 38844 11036
rect 38896 11024 38902 11076
rect 41785 11067 41843 11073
rect 41785 11033 41797 11067
rect 41831 11064 41843 11067
rect 54496 11064 54524 11104
rect 54570 11092 54576 11144
rect 54628 11132 54634 11144
rect 54628 11104 54673 11132
rect 54628 11092 54634 11104
rect 56226 11064 56232 11076
rect 41831 11036 45048 11064
rect 54496 11036 56232 11064
rect 41831 11033 41843 11036
rect 41785 11027 41843 11033
rect 37660 10968 37872 10996
rect 43530 10956 43536 11008
rect 43588 10996 43594 11008
rect 43806 10996 43812 11008
rect 43588 10968 43812 10996
rect 43588 10956 43594 10968
rect 43806 10956 43812 10968
rect 43864 10956 43870 11008
rect 45020 10996 45048 11036
rect 56226 11024 56232 11036
rect 56284 11024 56290 11076
rect 46385 10999 46443 11005
rect 46385 10996 46397 10999
rect 45020 10968 46397 10996
rect 46385 10965 46397 10968
rect 46431 10996 46443 10999
rect 46566 10996 46572 11008
rect 46431 10968 46572 10996
rect 46431 10965 46443 10968
rect 46385 10959 46443 10965
rect 46566 10956 46572 10968
rect 46624 10996 46630 11008
rect 46934 10996 46940 11008
rect 46624 10968 46940 10996
rect 46624 10956 46630 10968
rect 46934 10956 46940 10968
rect 46992 10956 46998 11008
rect 48406 10956 48412 11008
rect 48464 10996 48470 11008
rect 54570 10996 54576 11008
rect 48464 10968 54576 10996
rect 48464 10956 48470 10968
rect 54570 10956 54576 10968
rect 54628 10956 54634 11008
rect 56428 10996 56456 11163
rect 56686 11160 56692 11172
rect 56744 11160 56750 11212
rect 58897 11203 58955 11209
rect 58897 11169 58909 11203
rect 58943 11169 58955 11203
rect 58897 11163 58955 11169
rect 56594 11092 56600 11144
rect 56652 11132 56658 11144
rect 58912 11132 58940 11163
rect 56652 11104 58940 11132
rect 56652 11092 56658 11104
rect 57330 10996 57336 11008
rect 56428 10968 57336 10996
rect 57330 10956 57336 10968
rect 57388 10956 57394 11008
rect 1104 10906 62192 10928
rect 1104 10854 11163 10906
rect 11215 10854 11227 10906
rect 11279 10854 11291 10906
rect 11343 10854 11355 10906
rect 11407 10854 31526 10906
rect 31578 10854 31590 10906
rect 31642 10854 31654 10906
rect 31706 10854 31718 10906
rect 31770 10854 51888 10906
rect 51940 10854 51952 10906
rect 52004 10854 52016 10906
rect 52068 10854 52080 10906
rect 52132 10854 62192 10906
rect 1104 10832 62192 10854
rect 3142 10752 3148 10804
rect 3200 10792 3206 10804
rect 6638 10792 6644 10804
rect 3200 10764 6644 10792
rect 3200 10752 3206 10764
rect 6638 10752 6644 10764
rect 6696 10792 6702 10804
rect 7098 10792 7104 10804
rect 6696 10764 6868 10792
rect 7059 10764 7104 10792
rect 6696 10752 6702 10764
rect 3237 10659 3295 10665
rect 3237 10625 3249 10659
rect 3283 10656 3295 10659
rect 5442 10656 5448 10668
rect 3283 10628 5448 10656
rect 3283 10625 3295 10628
rect 3237 10619 3295 10625
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 6840 10656 6868 10764
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 7558 10752 7564 10804
rect 7616 10792 7622 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 7616 10764 8953 10792
rect 7616 10752 7622 10764
rect 8941 10761 8953 10764
rect 8987 10792 8999 10795
rect 9674 10792 9680 10804
rect 8987 10764 9680 10792
rect 8987 10761 8999 10764
rect 8941 10755 8999 10761
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 18414 10752 18420 10804
rect 18472 10792 18478 10804
rect 18785 10795 18843 10801
rect 18785 10792 18797 10795
rect 18472 10764 18797 10792
rect 18472 10752 18478 10764
rect 18785 10761 18797 10764
rect 18831 10761 18843 10795
rect 18785 10755 18843 10761
rect 14093 10727 14151 10733
rect 14093 10693 14105 10727
rect 14139 10724 14151 10727
rect 15010 10724 15016 10736
rect 14139 10696 15016 10724
rect 14139 10693 14151 10696
rect 14093 10687 14151 10693
rect 15010 10684 15016 10696
rect 15068 10684 15074 10736
rect 16390 10724 16396 10736
rect 16351 10696 16396 10724
rect 16390 10684 16396 10696
rect 16448 10724 16454 10736
rect 16666 10724 16672 10736
rect 16448 10696 16672 10724
rect 16448 10684 16454 10696
rect 16666 10684 16672 10696
rect 16724 10684 16730 10736
rect 6840 10628 11100 10656
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 2869 10591 2927 10597
rect 2869 10588 2881 10591
rect 2832 10560 2881 10588
rect 2832 10548 2838 10560
rect 2869 10557 2881 10560
rect 2915 10557 2927 10591
rect 2869 10551 2927 10557
rect 3970 10548 3976 10600
rect 4028 10588 4034 10600
rect 4065 10591 4123 10597
rect 4065 10588 4077 10591
rect 4028 10560 4077 10588
rect 4028 10548 4034 10560
rect 4065 10557 4077 10560
rect 4111 10557 4123 10591
rect 4065 10551 4123 10557
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10588 4399 10591
rect 6730 10588 6736 10600
rect 4387 10560 6736 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 6730 10548 6736 10560
rect 6788 10548 6794 10600
rect 6932 10597 6960 10628
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 6917 10591 6975 10597
rect 6917 10557 6929 10591
rect 6963 10557 6975 10591
rect 8754 10588 8760 10600
rect 8715 10560 8760 10588
rect 6917 10551 6975 10557
rect 2685 10523 2743 10529
rect 2685 10489 2697 10523
rect 2731 10489 2743 10523
rect 6840 10520 6868 10551
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 9858 10588 9864 10600
rect 9819 10560 9864 10588
rect 9858 10548 9864 10560
rect 9916 10548 9922 10600
rect 10962 10588 10968 10600
rect 10923 10560 10968 10588
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 11072 10597 11100 10628
rect 12158 10616 12164 10668
rect 12216 10656 12222 10668
rect 12529 10659 12587 10665
rect 12529 10656 12541 10659
rect 12216 10628 12541 10656
rect 12216 10616 12222 10628
rect 12529 10625 12541 10628
rect 12575 10625 12587 10659
rect 12529 10619 12587 10625
rect 12805 10659 12863 10665
rect 12805 10625 12817 10659
rect 12851 10656 12863 10659
rect 14458 10656 14464 10668
rect 12851 10628 14464 10656
rect 12851 10625 12863 10628
rect 12805 10619 12863 10625
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 18800 10656 18828 10755
rect 20898 10752 20904 10804
rect 20956 10792 20962 10804
rect 32306 10792 32312 10804
rect 20956 10764 32312 10792
rect 20956 10752 20962 10764
rect 32306 10752 32312 10764
rect 32364 10752 32370 10804
rect 33244 10764 34100 10792
rect 19061 10727 19119 10733
rect 19061 10693 19073 10727
rect 19107 10724 19119 10727
rect 20622 10724 20628 10736
rect 19107 10696 20628 10724
rect 19107 10693 19119 10696
rect 19061 10687 19119 10693
rect 20622 10684 20628 10696
rect 20680 10684 20686 10736
rect 33244 10733 33272 10764
rect 33229 10727 33287 10733
rect 33229 10693 33241 10727
rect 33275 10693 33287 10727
rect 33870 10724 33876 10736
rect 33229 10687 33287 10693
rect 33612 10696 33876 10724
rect 18800 10628 19564 10656
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10588 11115 10591
rect 11606 10588 11612 10600
rect 11103 10560 11612 10588
rect 11103 10557 11115 10560
rect 11057 10551 11115 10557
rect 11606 10548 11612 10560
rect 11664 10548 11670 10600
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10557 15071 10591
rect 15286 10588 15292 10600
rect 15247 10560 15292 10588
rect 15013 10551 15071 10557
rect 2685 10483 2743 10489
rect 5000 10492 6868 10520
rect 11517 10523 11575 10529
rect 2700 10452 2728 10483
rect 4062 10452 4068 10464
rect 2700 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10452 4126 10464
rect 5000 10452 5028 10492
rect 11517 10489 11529 10523
rect 11563 10520 11575 10523
rect 12066 10520 12072 10532
rect 11563 10492 12072 10520
rect 11563 10489 11575 10492
rect 11517 10483 11575 10489
rect 12066 10480 12072 10492
rect 12124 10480 12130 10532
rect 4120 10424 5028 10452
rect 5629 10455 5687 10461
rect 4120 10412 4126 10424
rect 5629 10421 5641 10455
rect 5675 10452 5687 10455
rect 7282 10452 7288 10464
rect 5675 10424 7288 10452
rect 5675 10421 5687 10424
rect 5629 10415 5687 10421
rect 7282 10412 7288 10424
rect 7340 10452 7346 10464
rect 7650 10452 7656 10464
rect 7340 10424 7656 10452
rect 7340 10412 7346 10424
rect 7650 10412 7656 10424
rect 7708 10412 7714 10464
rect 10042 10452 10048 10464
rect 10003 10424 10048 10452
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 10962 10412 10968 10464
rect 11020 10452 11026 10464
rect 13170 10452 13176 10464
rect 11020 10424 13176 10452
rect 11020 10412 11026 10424
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 15028 10452 15056 10551
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 16298 10548 16304 10600
rect 16356 10588 16362 10600
rect 18969 10591 19027 10597
rect 18969 10588 18981 10591
rect 16356 10560 18981 10588
rect 16356 10548 16362 10560
rect 18969 10557 18981 10560
rect 19015 10557 19027 10591
rect 18969 10551 19027 10557
rect 19334 10548 19340 10600
rect 19392 10588 19398 10600
rect 19536 10588 19564 10628
rect 19610 10616 19616 10668
rect 19668 10656 19674 10668
rect 19797 10659 19855 10665
rect 19797 10656 19809 10659
rect 19668 10628 19809 10656
rect 19668 10616 19674 10628
rect 19797 10625 19809 10628
rect 19843 10625 19855 10659
rect 21085 10659 21143 10665
rect 21085 10656 21097 10659
rect 19797 10619 19855 10625
rect 20640 10628 21097 10656
rect 19702 10588 19708 10600
rect 19392 10560 19437 10588
rect 19536 10560 19708 10588
rect 19392 10548 19398 10560
rect 19702 10548 19708 10560
rect 19760 10588 19766 10600
rect 20640 10588 20668 10628
rect 21085 10625 21097 10628
rect 21131 10656 21143 10659
rect 22186 10656 22192 10668
rect 21131 10628 22192 10656
rect 21131 10625 21143 10628
rect 21085 10619 21143 10625
rect 22186 10616 22192 10628
rect 22244 10616 22250 10668
rect 22741 10659 22799 10665
rect 22741 10625 22753 10659
rect 22787 10656 22799 10659
rect 24210 10656 24216 10668
rect 22787 10628 24216 10656
rect 22787 10625 22799 10628
rect 22741 10619 22799 10625
rect 24210 10616 24216 10628
rect 24268 10616 24274 10668
rect 24762 10616 24768 10668
rect 24820 10656 24826 10668
rect 25225 10659 25283 10665
rect 25225 10656 25237 10659
rect 24820 10628 25237 10656
rect 24820 10616 24826 10628
rect 25225 10625 25237 10628
rect 25271 10625 25283 10659
rect 25225 10619 25283 10625
rect 25866 10616 25872 10668
rect 25924 10656 25930 10668
rect 26605 10659 26663 10665
rect 26605 10656 26617 10659
rect 25924 10628 26617 10656
rect 25924 10616 25930 10628
rect 26605 10625 26617 10628
rect 26651 10625 26663 10659
rect 26605 10619 26663 10625
rect 26881 10659 26939 10665
rect 26881 10625 26893 10659
rect 26927 10656 26939 10659
rect 27062 10656 27068 10668
rect 26927 10628 27068 10656
rect 26927 10625 26939 10628
rect 26881 10619 26939 10625
rect 27062 10616 27068 10628
rect 27120 10616 27126 10668
rect 27614 10616 27620 10668
rect 27672 10656 27678 10668
rect 29733 10659 29791 10665
rect 29733 10656 29745 10659
rect 27672 10628 29745 10656
rect 27672 10616 27678 10628
rect 29733 10625 29745 10628
rect 29779 10625 29791 10659
rect 29733 10619 29791 10625
rect 20806 10588 20812 10600
rect 19760 10560 20668 10588
rect 20767 10560 20812 10588
rect 19760 10548 19766 10560
rect 20806 10548 20812 10560
rect 20864 10548 20870 10600
rect 21361 10591 21419 10597
rect 21361 10557 21373 10591
rect 21407 10588 21419 10591
rect 23566 10588 23572 10600
rect 21407 10560 23572 10588
rect 21407 10557 21419 10560
rect 21361 10551 21419 10557
rect 23566 10548 23572 10560
rect 23624 10548 23630 10600
rect 23661 10591 23719 10597
rect 23661 10557 23673 10591
rect 23707 10588 23719 10591
rect 25317 10591 25375 10597
rect 23707 10560 23980 10588
rect 23707 10557 23719 10560
rect 23661 10551 23719 10557
rect 19242 10520 19248 10532
rect 19203 10492 19248 10520
rect 19242 10480 19248 10492
rect 19300 10480 19306 10532
rect 19352 10492 20668 10520
rect 15746 10452 15752 10464
rect 15028 10424 15752 10452
rect 15746 10412 15752 10424
rect 15804 10412 15810 10464
rect 16390 10412 16396 10464
rect 16448 10452 16454 10464
rect 18966 10452 18972 10464
rect 16448 10424 18972 10452
rect 16448 10412 16454 10424
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 19058 10412 19064 10464
rect 19116 10452 19122 10464
rect 19352 10452 19380 10492
rect 19116 10424 19380 10452
rect 19116 10412 19122 10424
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 20162 10452 20168 10464
rect 19484 10424 20168 10452
rect 19484 10412 19490 10424
rect 20162 10412 20168 10424
rect 20220 10412 20226 10464
rect 20640 10461 20668 10492
rect 22554 10480 22560 10532
rect 22612 10520 22618 10532
rect 23676 10520 23704 10551
rect 22612 10492 23704 10520
rect 22612 10480 22618 10492
rect 20625 10455 20683 10461
rect 20625 10421 20637 10455
rect 20671 10421 20683 10455
rect 23842 10452 23848 10464
rect 23803 10424 23848 10452
rect 20625 10415 20683 10421
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 23952 10452 23980 10560
rect 25317 10557 25329 10591
rect 25363 10588 25375 10591
rect 25406 10588 25412 10600
rect 25363 10560 25412 10588
rect 25363 10557 25375 10560
rect 25317 10551 25375 10557
rect 25406 10548 25412 10560
rect 25464 10588 25470 10600
rect 28261 10591 28319 10597
rect 28261 10588 28273 10591
rect 25464 10560 28273 10588
rect 25464 10548 25470 10560
rect 28261 10557 28273 10560
rect 28307 10557 28319 10591
rect 28261 10551 28319 10557
rect 29457 10591 29515 10597
rect 29457 10557 29469 10591
rect 29503 10588 29515 10591
rect 30098 10588 30104 10600
rect 29503 10560 30104 10588
rect 29503 10557 29515 10560
rect 29457 10551 29515 10557
rect 30098 10548 30104 10560
rect 30156 10548 30162 10600
rect 30650 10588 30656 10600
rect 30611 10560 30656 10588
rect 30650 10548 30656 10560
rect 30708 10548 30714 10600
rect 31846 10588 31852 10600
rect 31807 10560 31852 10588
rect 31846 10548 31852 10560
rect 31904 10548 31910 10600
rect 33134 10548 33140 10600
rect 33192 10588 33198 10600
rect 33612 10597 33640 10696
rect 33870 10684 33876 10696
rect 33928 10684 33934 10736
rect 34072 10656 34100 10764
rect 36078 10752 36084 10804
rect 36136 10792 36142 10804
rect 36265 10795 36323 10801
rect 36265 10792 36277 10795
rect 36136 10764 36277 10792
rect 36136 10752 36142 10764
rect 36265 10761 36277 10764
rect 36311 10761 36323 10795
rect 43714 10792 43720 10804
rect 43675 10764 43720 10792
rect 36265 10755 36323 10761
rect 43714 10752 43720 10764
rect 43772 10752 43778 10804
rect 49050 10792 49056 10804
rect 48332 10764 49056 10792
rect 38473 10727 38531 10733
rect 38473 10693 38485 10727
rect 38519 10724 38531 10727
rect 39022 10724 39028 10736
rect 38519 10696 39028 10724
rect 38519 10693 38531 10696
rect 38473 10687 38531 10693
rect 39022 10684 39028 10696
rect 39080 10684 39086 10736
rect 35161 10659 35219 10665
rect 35161 10656 35173 10659
rect 34072 10628 35173 10656
rect 35161 10625 35173 10628
rect 35207 10625 35219 10659
rect 35161 10619 35219 10625
rect 39206 10616 39212 10668
rect 39264 10656 39270 10668
rect 42153 10659 42211 10665
rect 42153 10656 42165 10659
rect 39264 10628 42165 10656
rect 39264 10616 39270 10628
rect 42153 10625 42165 10628
rect 42199 10656 42211 10659
rect 42334 10656 42340 10668
rect 42199 10628 42340 10656
rect 42199 10625 42211 10628
rect 42153 10619 42211 10625
rect 42334 10616 42340 10628
rect 42392 10616 42398 10668
rect 45094 10656 45100 10668
rect 45055 10628 45100 10656
rect 45094 10616 45100 10628
rect 45152 10616 45158 10668
rect 46106 10656 46112 10668
rect 46067 10628 46112 10656
rect 46106 10616 46112 10628
rect 46164 10616 46170 10668
rect 48332 10665 48360 10764
rect 49050 10752 49056 10764
rect 49108 10752 49114 10804
rect 49881 10795 49939 10801
rect 49881 10761 49893 10795
rect 49927 10792 49939 10795
rect 50062 10792 50068 10804
rect 49927 10764 50068 10792
rect 49927 10761 49939 10764
rect 49881 10755 49939 10761
rect 50062 10752 50068 10764
rect 50120 10752 50126 10804
rect 53098 10752 53104 10804
rect 53156 10792 53162 10804
rect 53193 10795 53251 10801
rect 53193 10792 53205 10795
rect 53156 10764 53205 10792
rect 53156 10752 53162 10764
rect 53193 10761 53205 10764
rect 53239 10761 53251 10795
rect 53193 10755 53251 10761
rect 55677 10727 55735 10733
rect 55677 10693 55689 10727
rect 55723 10724 55735 10727
rect 56778 10724 56784 10736
rect 55723 10696 56784 10724
rect 55723 10693 55735 10696
rect 55677 10687 55735 10693
rect 56778 10684 56784 10696
rect 56836 10684 56842 10736
rect 48317 10659 48375 10665
rect 48317 10625 48329 10659
rect 48363 10625 48375 10659
rect 48317 10619 48375 10625
rect 52362 10616 52368 10668
rect 52420 10656 52426 10668
rect 57330 10656 57336 10668
rect 52420 10628 53052 10656
rect 57291 10628 57336 10656
rect 52420 10616 52426 10628
rect 33778 10597 33784 10600
rect 33413 10591 33471 10597
rect 33413 10588 33425 10591
rect 33192 10560 33425 10588
rect 33192 10548 33198 10560
rect 33413 10557 33425 10560
rect 33459 10557 33471 10591
rect 33413 10551 33471 10557
rect 33597 10591 33655 10597
rect 33597 10557 33609 10591
rect 33643 10557 33655 10591
rect 33597 10551 33655 10557
rect 33757 10591 33784 10597
rect 33757 10557 33769 10591
rect 33757 10551 33784 10557
rect 33778 10548 33784 10551
rect 33836 10548 33842 10600
rect 34882 10588 34888 10600
rect 34843 10560 34888 10588
rect 34882 10548 34888 10560
rect 34940 10548 34946 10600
rect 38654 10588 38660 10600
rect 38615 10560 38660 10588
rect 38654 10548 38660 10560
rect 38712 10548 38718 10600
rect 38838 10588 38844 10600
rect 38799 10560 38844 10588
rect 38838 10548 38844 10560
rect 38896 10548 38902 10600
rect 38930 10548 38936 10600
rect 38988 10588 38994 10600
rect 39025 10591 39083 10597
rect 39025 10588 39037 10591
rect 38988 10560 39037 10588
rect 38988 10548 38994 10560
rect 39025 10557 39037 10560
rect 39071 10557 39083 10591
rect 42426 10588 42432 10600
rect 42387 10560 42432 10588
rect 39025 10551 39083 10557
rect 42426 10548 42432 10560
rect 42484 10548 42490 10600
rect 44818 10588 44824 10600
rect 44779 10560 44824 10588
rect 44818 10548 44824 10560
rect 44876 10548 44882 10600
rect 45922 10548 45928 10600
rect 45980 10588 45986 10600
rect 46569 10591 46627 10597
rect 46569 10588 46581 10591
rect 45980 10560 46581 10588
rect 45980 10548 45986 10560
rect 46569 10557 46581 10560
rect 46615 10557 46627 10591
rect 46934 10588 46940 10600
rect 46895 10560 46940 10588
rect 46569 10551 46627 10557
rect 46934 10548 46940 10560
rect 46992 10548 46998 10600
rect 47029 10591 47087 10597
rect 47029 10557 47041 10591
rect 47075 10588 47087 10591
rect 47210 10588 47216 10600
rect 47075 10560 47216 10588
rect 47075 10557 47087 10560
rect 47029 10551 47087 10557
rect 47210 10548 47216 10560
rect 47268 10548 47274 10600
rect 48593 10591 48651 10597
rect 48593 10557 48605 10591
rect 48639 10588 48651 10591
rect 48958 10588 48964 10600
rect 48639 10560 48964 10588
rect 48639 10557 48651 10560
rect 48593 10551 48651 10557
rect 48958 10548 48964 10560
rect 49016 10548 49022 10600
rect 51721 10591 51779 10597
rect 51721 10588 51733 10591
rect 49252 10560 51733 10588
rect 25774 10520 25780 10532
rect 25735 10492 25780 10520
rect 25774 10480 25780 10492
rect 25832 10480 25838 10532
rect 27614 10480 27620 10532
rect 27672 10520 27678 10532
rect 29273 10523 29331 10529
rect 29273 10520 29285 10523
rect 27672 10492 29285 10520
rect 27672 10480 27678 10492
rect 29273 10489 29285 10492
rect 29319 10520 29331 10523
rect 30466 10520 30472 10532
rect 29319 10492 30472 10520
rect 29319 10489 29331 10492
rect 29273 10483 29331 10489
rect 30466 10480 30472 10492
rect 30524 10480 30530 10532
rect 44637 10523 44695 10529
rect 44637 10489 44649 10523
rect 44683 10520 44695 10523
rect 48406 10520 48412 10532
rect 44683 10492 48412 10520
rect 44683 10489 44695 10492
rect 44637 10483 44695 10489
rect 48406 10480 48412 10492
rect 48464 10480 48470 10532
rect 26142 10452 26148 10464
rect 23952 10424 26148 10452
rect 26142 10412 26148 10424
rect 26200 10412 26206 10464
rect 26878 10412 26884 10464
rect 26936 10452 26942 10464
rect 27522 10452 27528 10464
rect 26936 10424 27528 10452
rect 26936 10412 26942 10424
rect 27522 10412 27528 10424
rect 27580 10412 27586 10464
rect 30834 10452 30840 10464
rect 30795 10424 30840 10452
rect 30834 10412 30840 10424
rect 30892 10412 30898 10464
rect 32030 10452 32036 10464
rect 31991 10424 32036 10452
rect 32030 10412 32036 10424
rect 32088 10412 32094 10464
rect 46382 10412 46388 10464
rect 46440 10452 46446 10464
rect 49252 10452 49280 10560
rect 51721 10557 51733 10560
rect 51767 10557 51779 10591
rect 52914 10588 52920 10600
rect 52875 10560 52920 10588
rect 51721 10551 51779 10557
rect 49326 10480 49332 10532
rect 49384 10520 49390 10532
rect 51350 10520 51356 10532
rect 49384 10492 51356 10520
rect 49384 10480 49390 10492
rect 51350 10480 51356 10492
rect 51408 10480 51414 10532
rect 51736 10520 51764 10551
rect 52914 10548 52920 10560
rect 52972 10548 52978 10600
rect 53024 10597 53052 10628
rect 57330 10616 57336 10628
rect 57388 10616 57394 10668
rect 53009 10591 53067 10597
rect 53009 10557 53021 10591
rect 53055 10557 53067 10591
rect 54294 10588 54300 10600
rect 54255 10560 54300 10588
rect 53009 10551 53067 10557
rect 54294 10548 54300 10560
rect 54352 10548 54358 10600
rect 55398 10548 55404 10600
rect 55456 10588 55462 10600
rect 55861 10591 55919 10597
rect 55861 10588 55873 10591
rect 55456 10560 55873 10588
rect 55456 10548 55462 10560
rect 55861 10557 55873 10560
rect 55907 10557 55919 10591
rect 56042 10588 56048 10600
rect 56003 10560 56048 10588
rect 55861 10551 55919 10557
rect 56042 10548 56048 10560
rect 56100 10548 56106 10600
rect 56226 10588 56232 10600
rect 56187 10560 56232 10588
rect 56226 10548 56232 10560
rect 56284 10548 56290 10600
rect 57609 10591 57667 10597
rect 57609 10588 57621 10591
rect 57256 10560 57621 10588
rect 53190 10520 53196 10532
rect 51736 10492 53196 10520
rect 53190 10480 53196 10492
rect 53248 10480 53254 10532
rect 55766 10480 55772 10532
rect 55824 10520 55830 10532
rect 57256 10520 57284 10560
rect 57609 10557 57621 10560
rect 57655 10557 57667 10591
rect 57609 10551 57667 10557
rect 55824 10492 57284 10520
rect 55824 10480 55830 10492
rect 46440 10424 49280 10452
rect 46440 10412 46446 10424
rect 51442 10412 51448 10464
rect 51500 10452 51506 10464
rect 51813 10455 51871 10461
rect 51813 10452 51825 10455
rect 51500 10424 51825 10452
rect 51500 10412 51506 10424
rect 51813 10421 51825 10424
rect 51859 10421 51871 10455
rect 51813 10415 51871 10421
rect 54481 10455 54539 10461
rect 54481 10421 54493 10455
rect 54527 10452 54539 10455
rect 54754 10452 54760 10464
rect 54527 10424 54760 10452
rect 54527 10421 54539 10424
rect 54481 10415 54539 10421
rect 54754 10412 54760 10424
rect 54812 10412 54818 10464
rect 58710 10452 58716 10464
rect 58671 10424 58716 10452
rect 58710 10412 58716 10424
rect 58768 10412 58774 10464
rect 1104 10362 62192 10384
rect 1104 10310 21344 10362
rect 21396 10310 21408 10362
rect 21460 10310 21472 10362
rect 21524 10310 21536 10362
rect 21588 10310 41707 10362
rect 41759 10310 41771 10362
rect 41823 10310 41835 10362
rect 41887 10310 41899 10362
rect 41951 10310 62192 10362
rect 1104 10288 62192 10310
rect 5074 10208 5080 10260
rect 5132 10248 5138 10260
rect 5629 10251 5687 10257
rect 5629 10248 5641 10251
rect 5132 10220 5641 10248
rect 5132 10208 5138 10220
rect 5629 10217 5641 10220
rect 5675 10248 5687 10251
rect 10778 10248 10784 10260
rect 5675 10220 10784 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 11790 10208 11796 10260
rect 11848 10248 11854 10260
rect 12250 10248 12256 10260
rect 11848 10220 12256 10248
rect 11848 10208 11854 10220
rect 12250 10208 12256 10220
rect 12308 10248 12314 10260
rect 12308 10220 15976 10248
rect 12308 10208 12314 10220
rect 7006 10140 7012 10192
rect 7064 10180 7070 10192
rect 7101 10183 7159 10189
rect 7101 10180 7113 10183
rect 7064 10152 7113 10180
rect 7064 10140 7070 10152
rect 7101 10149 7113 10152
rect 7147 10149 7159 10183
rect 7101 10143 7159 10149
rect 11425 10183 11483 10189
rect 11425 10149 11437 10183
rect 11471 10180 11483 10183
rect 13722 10180 13728 10192
rect 11471 10152 13728 10180
rect 11471 10149 11483 10152
rect 11425 10143 11483 10149
rect 13722 10140 13728 10152
rect 13780 10140 13786 10192
rect 15102 10140 15108 10192
rect 15160 10180 15166 10192
rect 15289 10183 15347 10189
rect 15289 10180 15301 10183
rect 15160 10152 15301 10180
rect 15160 10140 15166 10152
rect 15289 10149 15301 10152
rect 15335 10149 15347 10183
rect 15289 10143 15347 10149
rect 15378 10140 15384 10192
rect 15436 10180 15442 10192
rect 15948 10180 15976 10220
rect 19242 10208 19248 10260
rect 19300 10248 19306 10260
rect 29730 10248 29736 10260
rect 19300 10220 29736 10248
rect 19300 10208 19306 10220
rect 29730 10208 29736 10220
rect 29788 10208 29794 10260
rect 34974 10248 34980 10260
rect 34935 10220 34980 10248
rect 34974 10208 34980 10220
rect 35032 10208 35038 10260
rect 36354 10248 36360 10260
rect 36315 10220 36360 10248
rect 36354 10208 36360 10220
rect 36412 10208 36418 10260
rect 38764 10220 44220 10248
rect 19521 10183 19579 10189
rect 19521 10180 19533 10183
rect 15436 10152 15884 10180
rect 15948 10152 19533 10180
rect 15436 10140 15442 10152
rect 15856 10124 15884 10152
rect 19521 10149 19533 10152
rect 19567 10149 19579 10183
rect 19521 10143 19579 10149
rect 19610 10140 19616 10192
rect 19668 10180 19674 10192
rect 23845 10183 23903 10189
rect 19668 10152 19713 10180
rect 19668 10140 19674 10152
rect 23845 10149 23857 10183
rect 23891 10180 23903 10183
rect 24762 10180 24768 10192
rect 23891 10152 24768 10180
rect 23891 10149 23903 10152
rect 23845 10143 23903 10149
rect 24762 10140 24768 10152
rect 24820 10140 24826 10192
rect 25593 10183 25651 10189
rect 25593 10180 25605 10183
rect 24872 10152 25605 10180
rect 6638 10112 6644 10124
rect 6599 10084 6644 10112
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 10042 10112 10048 10124
rect 9955 10084 10048 10112
rect 10042 10072 10048 10084
rect 10100 10112 10106 10124
rect 11606 10112 11612 10124
rect 10100 10084 11612 10112
rect 10100 10072 10106 10084
rect 11606 10072 11612 10084
rect 11664 10112 11670 10124
rect 11882 10112 11888 10124
rect 11664 10084 11888 10112
rect 11664 10072 11670 10084
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 12066 10112 12072 10124
rect 12027 10084 12072 10112
rect 12066 10072 12072 10084
rect 12124 10072 12130 10124
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10081 12495 10115
rect 12437 10075 12495 10081
rect 12621 10115 12679 10121
rect 12621 10081 12633 10115
rect 12667 10112 12679 10115
rect 13354 10112 13360 10124
rect 12667 10084 13360 10112
rect 12667 10081 12679 10084
rect 12621 10075 12679 10081
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 4028 10016 4077 10044
rect 4028 10004 4034 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4338 10044 4344 10056
rect 4299 10016 4344 10044
rect 4065 10007 4123 10013
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 6546 10044 6552 10056
rect 6507 10016 6552 10044
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 9953 10047 10011 10053
rect 9953 10044 9965 10047
rect 9732 10016 9965 10044
rect 9732 10004 9738 10016
rect 9953 10013 9965 10016
rect 9999 10013 10011 10047
rect 9953 10007 10011 10013
rect 10870 10004 10876 10056
rect 10928 10044 10934 10056
rect 11977 10047 12035 10053
rect 11977 10044 11989 10047
rect 10928 10016 11989 10044
rect 10928 10004 10934 10016
rect 11977 10013 11989 10016
rect 12023 10013 12035 10047
rect 12452 10044 12480 10075
rect 13354 10072 13360 10084
rect 13412 10072 13418 10124
rect 13449 10115 13507 10121
rect 13449 10081 13461 10115
rect 13495 10081 13507 10115
rect 13449 10075 13507 10081
rect 13170 10044 13176 10056
rect 12452 10016 13176 10044
rect 11977 10007 12035 10013
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 13464 9988 13492 10075
rect 15010 10072 15016 10124
rect 15068 10112 15074 10124
rect 15749 10115 15807 10121
rect 15749 10112 15761 10115
rect 15068 10084 15761 10112
rect 15068 10072 15074 10084
rect 15749 10081 15761 10084
rect 15795 10081 15807 10115
rect 15749 10075 15807 10081
rect 15838 10072 15844 10124
rect 15896 10112 15902 10124
rect 15933 10115 15991 10121
rect 15933 10112 15945 10115
rect 15896 10084 15945 10112
rect 15896 10072 15902 10084
rect 15933 10081 15945 10084
rect 15979 10081 15991 10115
rect 16114 10112 16120 10124
rect 16075 10084 16120 10112
rect 15933 10075 15991 10081
rect 16114 10072 16120 10084
rect 16172 10072 16178 10124
rect 17957 10115 18015 10121
rect 17957 10081 17969 10115
rect 18003 10112 18015 10115
rect 18414 10112 18420 10124
rect 18003 10084 18420 10112
rect 18003 10081 18015 10084
rect 17957 10075 18015 10081
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 19426 10112 19432 10124
rect 19387 10084 19432 10112
rect 19426 10072 19432 10084
rect 19484 10072 19490 10124
rect 21082 10112 21088 10124
rect 21043 10084 21088 10112
rect 21082 10072 21088 10084
rect 21140 10072 21146 10124
rect 21266 10072 21272 10124
rect 21324 10112 21330 10124
rect 21818 10112 21824 10124
rect 21324 10084 21824 10112
rect 21324 10072 21330 10084
rect 21818 10072 21824 10084
rect 21876 10112 21882 10124
rect 21876 10084 22140 10112
rect 21876 10072 21882 10084
rect 13814 10044 13820 10056
rect 13775 10016 13820 10044
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 17586 10004 17592 10056
rect 17644 10044 17650 10056
rect 17865 10047 17923 10053
rect 17865 10044 17877 10047
rect 17644 10016 17877 10044
rect 17644 10004 17650 10016
rect 17865 10013 17877 10016
rect 17911 10013 17923 10047
rect 17865 10007 17923 10013
rect 19245 10047 19303 10053
rect 19245 10013 19257 10047
rect 19291 10044 19303 10047
rect 19334 10044 19340 10056
rect 19291 10016 19340 10044
rect 19291 10013 19303 10016
rect 19245 10007 19303 10013
rect 19334 10004 19340 10016
rect 19392 10004 19398 10056
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10044 20039 10047
rect 22112 10044 22140 10084
rect 22186 10072 22192 10124
rect 22244 10112 22250 10124
rect 22465 10115 22523 10121
rect 22244 10084 22289 10112
rect 22244 10072 22250 10084
rect 22465 10081 22477 10115
rect 22511 10112 22523 10115
rect 23382 10112 23388 10124
rect 22511 10084 23388 10112
rect 22511 10081 22523 10084
rect 22465 10075 22523 10081
rect 23382 10072 23388 10084
rect 23440 10072 23446 10124
rect 23566 10072 23572 10124
rect 23624 10112 23630 10124
rect 24872 10112 24900 10152
rect 25593 10149 25605 10152
rect 25639 10149 25651 10183
rect 25593 10143 25651 10149
rect 25774 10140 25780 10192
rect 25832 10180 25838 10192
rect 28813 10183 28871 10189
rect 28813 10180 28825 10183
rect 25832 10152 28825 10180
rect 25832 10140 25838 10152
rect 28813 10149 28825 10152
rect 28859 10149 28871 10183
rect 28813 10143 28871 10149
rect 36081 10183 36139 10189
rect 36081 10149 36093 10183
rect 36127 10180 36139 10183
rect 38764 10180 38792 10220
rect 36127 10152 38792 10180
rect 39393 10183 39451 10189
rect 36127 10149 36139 10152
rect 36081 10143 36139 10149
rect 39393 10149 39405 10183
rect 39439 10180 39451 10183
rect 39482 10180 39488 10192
rect 39439 10152 39488 10180
rect 39439 10149 39451 10152
rect 39393 10143 39451 10149
rect 39482 10140 39488 10152
rect 39540 10140 39546 10192
rect 41414 10140 41420 10192
rect 41472 10180 41478 10192
rect 43714 10180 43720 10192
rect 41472 10152 43720 10180
rect 41472 10140 41478 10152
rect 25038 10112 25044 10124
rect 23624 10084 24900 10112
rect 24999 10084 25044 10112
rect 23624 10072 23630 10084
rect 25038 10072 25044 10084
rect 25096 10072 25102 10124
rect 25133 10115 25191 10121
rect 25133 10081 25145 10115
rect 25179 10112 25191 10115
rect 26418 10112 26424 10124
rect 25179 10084 26424 10112
rect 25179 10081 25191 10084
rect 25133 10075 25191 10081
rect 26418 10072 26424 10084
rect 26476 10072 26482 10124
rect 26789 10115 26847 10121
rect 26789 10081 26801 10115
rect 26835 10112 26847 10115
rect 26878 10112 26884 10124
rect 26835 10084 26884 10112
rect 26835 10081 26847 10084
rect 26789 10075 26847 10081
rect 26878 10072 26884 10084
rect 26936 10072 26942 10124
rect 27062 10112 27068 10124
rect 27023 10084 27068 10112
rect 27062 10072 27068 10084
rect 27120 10072 27126 10124
rect 27525 10115 27583 10121
rect 27525 10081 27537 10115
rect 27571 10112 27583 10115
rect 27614 10112 27620 10124
rect 27571 10084 27620 10112
rect 27571 10081 27583 10084
rect 27525 10075 27583 10081
rect 27614 10072 27620 10084
rect 27672 10072 27678 10124
rect 27709 10115 27767 10121
rect 27709 10081 27721 10115
rect 27755 10081 27767 10115
rect 28994 10112 29000 10124
rect 28955 10084 29000 10112
rect 27709 10075 27767 10081
rect 24670 10044 24676 10056
rect 20027 10016 22048 10044
rect 22112 10016 24676 10044
rect 20027 10013 20039 10016
rect 19981 10007 20039 10013
rect 11698 9936 11704 9988
rect 11756 9976 11762 9988
rect 12066 9976 12072 9988
rect 11756 9948 12072 9976
rect 11756 9936 11762 9948
rect 12066 9936 12072 9948
rect 12124 9936 12130 9988
rect 13446 9976 13452 9988
rect 13359 9948 13452 9976
rect 13446 9936 13452 9948
rect 13504 9976 13510 9988
rect 19610 9976 19616 9988
rect 13504 9948 19616 9976
rect 13504 9936 13510 9948
rect 19610 9936 19616 9948
rect 19668 9936 19674 9988
rect 21266 9976 21272 9988
rect 21227 9948 21272 9976
rect 21266 9936 21272 9948
rect 21324 9936 21330 9988
rect 10226 9908 10232 9920
rect 10187 9880 10232 9908
rect 10226 9868 10232 9880
rect 10284 9868 10290 9920
rect 11514 9868 11520 9920
rect 11572 9908 11578 9920
rect 13587 9911 13645 9917
rect 13587 9908 13599 9911
rect 11572 9880 13599 9908
rect 11572 9868 11578 9880
rect 13587 9877 13599 9880
rect 13633 9877 13645 9911
rect 13722 9908 13728 9920
rect 13683 9880 13728 9908
rect 13587 9871 13645 9877
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 14093 9911 14151 9917
rect 14093 9877 14105 9911
rect 14139 9908 14151 9911
rect 16022 9908 16028 9920
rect 14139 9880 16028 9908
rect 14139 9877 14151 9880
rect 14093 9871 14151 9877
rect 16022 9868 16028 9880
rect 16080 9868 16086 9920
rect 18141 9911 18199 9917
rect 18141 9877 18153 9911
rect 18187 9908 18199 9911
rect 21174 9908 21180 9920
rect 18187 9880 21180 9908
rect 18187 9877 18199 9880
rect 18141 9871 18199 9877
rect 21174 9868 21180 9880
rect 21232 9868 21238 9920
rect 22020 9908 22048 10016
rect 24670 10004 24676 10016
rect 24728 10004 24734 10056
rect 25314 10004 25320 10056
rect 25372 10044 25378 10056
rect 27724 10044 27752 10075
rect 28994 10072 29000 10084
rect 29052 10072 29058 10124
rect 30193 10115 30251 10121
rect 30193 10081 30205 10115
rect 30239 10112 30251 10115
rect 30650 10112 30656 10124
rect 30239 10084 30656 10112
rect 30239 10081 30251 10084
rect 30193 10075 30251 10081
rect 30650 10072 30656 10084
rect 30708 10112 30714 10124
rect 32122 10112 32128 10124
rect 30708 10084 32128 10112
rect 30708 10072 30714 10084
rect 32122 10072 32128 10084
rect 32180 10072 32186 10124
rect 32306 10112 32312 10124
rect 32267 10084 32312 10112
rect 32306 10072 32312 10084
rect 32364 10072 32370 10124
rect 33594 10112 33600 10124
rect 33555 10084 33600 10112
rect 33594 10072 33600 10084
rect 33652 10072 33658 10124
rect 34146 10072 34152 10124
rect 34204 10112 34210 10124
rect 36265 10115 36323 10121
rect 36265 10112 36277 10115
rect 34204 10084 36277 10112
rect 34204 10072 34210 10084
rect 36265 10081 36277 10084
rect 36311 10081 36323 10115
rect 37734 10112 37740 10124
rect 37695 10084 37740 10112
rect 36265 10075 36323 10081
rect 37734 10072 37740 10084
rect 37792 10072 37798 10124
rect 39574 10072 39580 10124
rect 39632 10112 39638 10124
rect 39853 10115 39911 10121
rect 39853 10112 39865 10115
rect 39632 10084 39865 10112
rect 39632 10072 39638 10084
rect 39853 10081 39865 10084
rect 39899 10081 39911 10115
rect 39853 10075 39911 10081
rect 40037 10115 40095 10121
rect 40037 10081 40049 10115
rect 40083 10081 40095 10115
rect 40037 10075 40095 10081
rect 40221 10115 40279 10121
rect 40221 10081 40233 10115
rect 40267 10112 40279 10115
rect 40494 10112 40500 10124
rect 40267 10084 40500 10112
rect 40267 10081 40279 10084
rect 40221 10075 40279 10081
rect 32214 10044 32220 10056
rect 25372 10016 27752 10044
rect 32175 10016 32220 10044
rect 25372 10004 25378 10016
rect 32214 10004 32220 10016
rect 32272 10004 32278 10056
rect 32769 10047 32827 10053
rect 32769 10013 32781 10047
rect 32815 10044 32827 10047
rect 33410 10044 33416 10056
rect 32815 10016 33416 10044
rect 32815 10013 32827 10016
rect 32769 10007 32827 10013
rect 33410 10004 33416 10016
rect 33468 10004 33474 10056
rect 33873 10047 33931 10053
rect 33873 10013 33885 10047
rect 33919 10044 33931 10047
rect 35618 10044 35624 10056
rect 33919 10016 35624 10044
rect 33919 10013 33931 10016
rect 33873 10007 33931 10013
rect 35618 10004 35624 10016
rect 35676 10004 35682 10056
rect 38838 10004 38844 10056
rect 38896 10044 38902 10056
rect 40052 10044 40080 10075
rect 40494 10072 40500 10084
rect 40552 10072 40558 10124
rect 41598 10072 41604 10124
rect 41656 10112 41662 10124
rect 42076 10121 42104 10152
rect 43714 10140 43720 10152
rect 43772 10140 43778 10192
rect 41693 10115 41751 10121
rect 41693 10112 41705 10115
rect 41656 10084 41705 10112
rect 41656 10072 41662 10084
rect 41693 10081 41705 10084
rect 41739 10081 41751 10115
rect 41693 10075 41751 10081
rect 42061 10115 42119 10121
rect 42061 10081 42073 10115
rect 42107 10081 42119 10115
rect 42061 10075 42119 10081
rect 42150 10072 42156 10124
rect 42208 10112 42214 10124
rect 42208 10084 42253 10112
rect 42208 10072 42214 10084
rect 42168 10044 42196 10072
rect 38896 10016 42196 10044
rect 38896 10004 38902 10016
rect 23290 9936 23296 9988
rect 23348 9976 23354 9988
rect 26605 9979 26663 9985
rect 26605 9976 26617 9979
rect 23348 9948 26617 9976
rect 23348 9936 23354 9948
rect 26605 9945 26617 9948
rect 26651 9945 26663 9979
rect 26605 9939 26663 9945
rect 26694 9936 26700 9988
rect 26752 9976 26758 9988
rect 27430 9976 27436 9988
rect 26752 9948 27436 9976
rect 26752 9936 26758 9948
rect 27430 9936 27436 9948
rect 27488 9936 27494 9988
rect 27706 9936 27712 9988
rect 27764 9976 27770 9988
rect 30377 9979 30435 9985
rect 30377 9976 30389 9979
rect 27764 9948 30389 9976
rect 27764 9936 27770 9948
rect 30377 9945 30389 9948
rect 30423 9945 30435 9979
rect 30377 9939 30435 9945
rect 41509 9979 41567 9985
rect 41509 9945 41521 9979
rect 41555 9976 41567 9979
rect 42426 9976 42432 9988
rect 41555 9948 42432 9976
rect 41555 9945 41567 9948
rect 41509 9939 41567 9945
rect 42426 9936 42432 9948
rect 42484 9936 42490 9988
rect 22922 9908 22928 9920
rect 22020 9880 22928 9908
rect 22922 9868 22928 9880
rect 22980 9868 22986 9920
rect 25038 9868 25044 9920
rect 25096 9908 25102 9920
rect 26712 9908 26740 9936
rect 25096 9880 26740 9908
rect 25096 9868 25102 9880
rect 27614 9868 27620 9920
rect 27672 9908 27678 9920
rect 29089 9911 29147 9917
rect 29089 9908 29101 9911
rect 27672 9880 29101 9908
rect 27672 9868 27678 9880
rect 29089 9877 29101 9880
rect 29135 9877 29147 9911
rect 29089 9871 29147 9877
rect 36906 9868 36912 9920
rect 36964 9908 36970 9920
rect 37921 9911 37979 9917
rect 37921 9908 37933 9911
rect 36964 9880 37933 9908
rect 36964 9868 36970 9880
rect 37921 9877 37933 9880
rect 37967 9877 37979 9911
rect 44192 9908 44220 10220
rect 44910 10208 44916 10260
rect 44968 10248 44974 10260
rect 47029 10251 47087 10257
rect 47029 10248 47041 10251
rect 44968 10220 47041 10248
rect 44968 10208 44974 10220
rect 47029 10217 47041 10220
rect 47075 10248 47087 10251
rect 47486 10248 47492 10260
rect 47075 10220 47492 10248
rect 47075 10217 47087 10220
rect 47029 10211 47087 10217
rect 47486 10208 47492 10220
rect 47544 10208 47550 10260
rect 49326 10248 49332 10260
rect 48792 10220 49332 10248
rect 47210 10140 47216 10192
rect 47268 10180 47274 10192
rect 48792 10180 48820 10220
rect 49326 10208 49332 10220
rect 49384 10208 49390 10260
rect 59354 10248 59360 10260
rect 56244 10220 59360 10248
rect 48958 10180 48964 10192
rect 47268 10152 48820 10180
rect 48919 10152 48964 10180
rect 47268 10140 47274 10152
rect 48958 10140 48964 10152
rect 49016 10140 49022 10192
rect 55766 10180 55772 10192
rect 55727 10152 55772 10180
rect 55766 10140 55772 10152
rect 55824 10140 55830 10192
rect 44361 10115 44419 10121
rect 44361 10081 44373 10115
rect 44407 10112 44419 10115
rect 45094 10112 45100 10124
rect 44407 10084 45100 10112
rect 44407 10081 44419 10084
rect 44361 10075 44419 10081
rect 45094 10072 45100 10084
rect 45152 10072 45158 10124
rect 46017 10115 46075 10121
rect 46017 10081 46029 10115
rect 46063 10112 46075 10115
rect 46106 10112 46112 10124
rect 46063 10084 46112 10112
rect 46063 10081 46075 10084
rect 46017 10075 46075 10081
rect 46106 10072 46112 10084
rect 46164 10112 46170 10124
rect 46845 10115 46903 10121
rect 46845 10112 46857 10115
rect 46164 10084 46857 10112
rect 46164 10072 46170 10084
rect 46845 10081 46857 10084
rect 46891 10081 46903 10115
rect 46845 10075 46903 10081
rect 49421 10115 49479 10121
rect 49421 10081 49433 10115
rect 49467 10112 49479 10115
rect 49510 10112 49516 10124
rect 49467 10084 49516 10112
rect 49467 10081 49479 10084
rect 49421 10075 49479 10081
rect 49510 10072 49516 10084
rect 49568 10072 49574 10124
rect 49789 10115 49847 10121
rect 49789 10081 49801 10115
rect 49835 10112 49847 10115
rect 50062 10112 50068 10124
rect 49835 10084 50068 10112
rect 49835 10081 49847 10084
rect 49789 10075 49847 10081
rect 50062 10072 50068 10084
rect 50120 10072 50126 10124
rect 51350 10072 51356 10124
rect 51408 10112 51414 10124
rect 54662 10112 54668 10124
rect 51408 10084 54524 10112
rect 54623 10084 54668 10112
rect 51408 10072 51414 10084
rect 44634 10044 44640 10056
rect 44595 10016 44640 10044
rect 44634 10004 44640 10016
rect 44692 10004 44698 10056
rect 49694 10004 49700 10056
rect 49752 10044 49758 10056
rect 49881 10047 49939 10053
rect 49881 10044 49893 10047
rect 49752 10016 49893 10044
rect 49752 10004 49758 10016
rect 49881 10013 49893 10016
rect 49927 10013 49939 10047
rect 51534 10044 51540 10056
rect 51495 10016 51540 10044
rect 49881 10007 49939 10013
rect 51534 10004 51540 10016
rect 51592 10004 51598 10056
rect 51718 10004 51724 10056
rect 51776 10044 51782 10056
rect 51813 10047 51871 10053
rect 51813 10044 51825 10047
rect 51776 10016 51825 10044
rect 51776 10004 51782 10016
rect 51813 10013 51825 10016
rect 51859 10013 51871 10047
rect 51813 10007 51871 10013
rect 54496 9976 54524 10084
rect 54662 10072 54668 10084
rect 54720 10072 54726 10124
rect 56244 10121 56272 10220
rect 59354 10208 59360 10220
rect 59412 10208 59418 10260
rect 56229 10115 56287 10121
rect 56229 10081 56241 10115
rect 56275 10081 56287 10115
rect 56229 10075 56287 10081
rect 56597 10115 56655 10121
rect 56597 10081 56609 10115
rect 56643 10112 56655 10115
rect 58710 10112 58716 10124
rect 56643 10084 58716 10112
rect 56643 10081 56655 10084
rect 56597 10075 56655 10081
rect 54570 10004 54576 10056
rect 54628 10044 54634 10056
rect 56612 10044 56640 10075
rect 58710 10072 58716 10084
rect 58768 10072 58774 10124
rect 54628 10016 56640 10044
rect 56689 10047 56747 10053
rect 54628 10004 54634 10016
rect 56689 10013 56701 10047
rect 56735 10013 56747 10047
rect 56689 10007 56747 10013
rect 56594 9976 56600 9988
rect 54496 9948 56600 9976
rect 56594 9936 56600 9948
rect 56652 9976 56658 9988
rect 56704 9976 56732 10007
rect 57330 10004 57336 10056
rect 57388 10044 57394 10056
rect 57609 10047 57667 10053
rect 57609 10044 57621 10047
rect 57388 10016 57621 10044
rect 57388 10004 57394 10016
rect 57609 10013 57621 10016
rect 57655 10013 57667 10047
rect 57609 10007 57667 10013
rect 57885 10047 57943 10053
rect 57885 10013 57897 10047
rect 57931 10044 57943 10047
rect 58066 10044 58072 10056
rect 57931 10016 58072 10044
rect 57931 10013 57943 10016
rect 57885 10007 57943 10013
rect 58066 10004 58072 10016
rect 58124 10004 58130 10056
rect 56652 9948 56732 9976
rect 56652 9936 56658 9948
rect 50246 9908 50252 9920
rect 44192 9880 50252 9908
rect 37921 9871 37979 9877
rect 50246 9868 50252 9880
rect 50304 9868 50310 9920
rect 53101 9911 53159 9917
rect 53101 9877 53113 9911
rect 53147 9908 53159 9911
rect 53190 9908 53196 9920
rect 53147 9880 53196 9908
rect 53147 9877 53159 9880
rect 53101 9871 53159 9877
rect 53190 9868 53196 9880
rect 53248 9868 53254 9920
rect 54846 9908 54852 9920
rect 54807 9880 54852 9908
rect 54846 9868 54852 9880
rect 54904 9868 54910 9920
rect 58526 9868 58532 9920
rect 58584 9908 58590 9920
rect 58989 9911 59047 9917
rect 58989 9908 59001 9911
rect 58584 9880 59001 9908
rect 58584 9868 58590 9880
rect 58989 9877 59001 9880
rect 59035 9877 59047 9911
rect 58989 9871 59047 9877
rect 1104 9818 62192 9840
rect 1104 9766 11163 9818
rect 11215 9766 11227 9818
rect 11279 9766 11291 9818
rect 11343 9766 11355 9818
rect 11407 9766 31526 9818
rect 31578 9766 31590 9818
rect 31642 9766 31654 9818
rect 31706 9766 31718 9818
rect 31770 9766 51888 9818
rect 51940 9766 51952 9818
rect 52004 9766 52016 9818
rect 52068 9766 52080 9818
rect 52132 9766 62192 9818
rect 1104 9744 62192 9766
rect 9858 9664 9864 9716
rect 9916 9704 9922 9716
rect 10229 9707 10287 9713
rect 10229 9704 10241 9707
rect 9916 9676 10241 9704
rect 9916 9664 9922 9676
rect 10229 9673 10241 9676
rect 10275 9704 10287 9707
rect 13446 9704 13452 9716
rect 10275 9676 13452 9704
rect 10275 9673 10287 9676
rect 10229 9667 10287 9673
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 37001 9707 37059 9713
rect 37001 9673 37013 9707
rect 37047 9673 37059 9707
rect 37001 9667 37059 9673
rect 6730 9596 6736 9648
rect 6788 9636 6794 9648
rect 7101 9639 7159 9645
rect 7101 9636 7113 9639
rect 6788 9608 7113 9636
rect 6788 9596 6794 9608
rect 7101 9605 7113 9608
rect 7147 9605 7159 9639
rect 7101 9599 7159 9605
rect 15197 9639 15255 9645
rect 15197 9605 15209 9639
rect 15243 9636 15255 9639
rect 15286 9636 15292 9648
rect 15243 9608 15292 9636
rect 15243 9605 15255 9608
rect 15197 9599 15255 9605
rect 15286 9596 15292 9608
rect 15344 9596 15350 9648
rect 17037 9639 17095 9645
rect 17037 9605 17049 9639
rect 17083 9636 17095 9639
rect 17494 9636 17500 9648
rect 17083 9608 17500 9636
rect 17083 9605 17095 9608
rect 17037 9599 17095 9605
rect 17494 9596 17500 9608
rect 17552 9596 17558 9648
rect 19610 9636 19616 9648
rect 17604 9608 19616 9636
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9568 3019 9571
rect 3970 9568 3976 9580
rect 3007 9540 3976 9568
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3970 9528 3976 9540
rect 4028 9528 4034 9580
rect 10962 9568 10968 9580
rect 4356 9540 10968 9568
rect 3234 9500 3240 9512
rect 3195 9472 3240 9500
rect 3234 9460 3240 9472
rect 3292 9460 3298 9512
rect 2958 9324 2964 9376
rect 3016 9364 3022 9376
rect 4356 9373 4384 9540
rect 10962 9528 10968 9540
rect 11020 9528 11026 9580
rect 12158 9528 12164 9580
rect 12216 9568 12222 9580
rect 12437 9571 12495 9577
rect 12437 9568 12449 9571
rect 12216 9540 12449 9568
rect 12216 9528 12222 9540
rect 12437 9537 12449 9540
rect 12483 9537 12495 9571
rect 15838 9568 15844 9580
rect 15799 9540 15844 9568
rect 12437 9531 12495 9537
rect 15838 9528 15844 9540
rect 15896 9528 15902 9580
rect 16666 9568 16672 9580
rect 16500 9540 16672 9568
rect 7190 9460 7196 9512
rect 7248 9500 7254 9512
rect 7285 9503 7343 9509
rect 7285 9500 7297 9503
rect 7248 9472 7297 9500
rect 7248 9460 7254 9472
rect 7285 9469 7297 9472
rect 7331 9469 7343 9503
rect 7466 9500 7472 9512
rect 7427 9472 7472 9500
rect 7285 9463 7343 9469
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 7650 9500 7656 9512
rect 7611 9472 7656 9500
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9500 8999 9503
rect 11054 9500 11060 9512
rect 8987 9472 11060 9500
rect 8987 9469 8999 9472
rect 8941 9463 8999 9469
rect 8680 9376 8708 9463
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9500 11207 9503
rect 11514 9500 11520 9512
rect 11195 9472 11520 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 11514 9460 11520 9472
rect 11572 9460 11578 9512
rect 12176 9432 12204 9528
rect 12710 9500 12716 9512
rect 12671 9472 12716 9500
rect 12710 9460 12716 9472
rect 12768 9460 12774 9512
rect 12986 9460 12992 9512
rect 13044 9500 13050 9512
rect 13722 9500 13728 9512
rect 13044 9472 13728 9500
rect 13044 9460 13050 9472
rect 13722 9460 13728 9472
rect 13780 9500 13786 9512
rect 15378 9500 15384 9512
rect 13780 9472 14780 9500
rect 15339 9472 15384 9500
rect 13780 9460 13786 9472
rect 9600 9404 12204 9432
rect 4341 9367 4399 9373
rect 4341 9364 4353 9367
rect 3016 9336 4353 9364
rect 3016 9324 3022 9336
rect 4341 9333 4353 9336
rect 4387 9333 4399 9367
rect 8662 9364 8668 9376
rect 8575 9336 8668 9364
rect 4341 9327 4399 9333
rect 8662 9324 8668 9336
rect 8720 9364 8726 9376
rect 9600 9364 9628 9404
rect 13814 9392 13820 9444
rect 13872 9432 13878 9444
rect 14093 9435 14151 9441
rect 14093 9432 14105 9435
rect 13872 9404 14105 9432
rect 13872 9392 13878 9404
rect 14093 9401 14105 9404
rect 14139 9432 14151 9435
rect 14642 9432 14648 9444
rect 14139 9404 14648 9432
rect 14139 9401 14151 9404
rect 14093 9395 14151 9401
rect 14642 9392 14648 9404
rect 14700 9392 14706 9444
rect 14752 9432 14780 9472
rect 15378 9460 15384 9472
rect 15436 9460 15442 9512
rect 15749 9503 15807 9509
rect 15749 9469 15761 9503
rect 15795 9500 15807 9503
rect 16500 9500 16528 9540
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 15795 9472 16528 9500
rect 15795 9469 15807 9472
rect 15749 9463 15807 9469
rect 16574 9460 16580 9512
rect 16632 9500 16638 9512
rect 16853 9503 16911 9509
rect 16853 9500 16865 9503
rect 16632 9472 16865 9500
rect 16632 9460 16638 9472
rect 16853 9469 16865 9472
rect 16899 9500 16911 9503
rect 17604 9500 17632 9608
rect 19610 9596 19616 9608
rect 19668 9596 19674 9648
rect 20714 9596 20720 9648
rect 20772 9636 20778 9648
rect 23106 9636 23112 9648
rect 20772 9608 23112 9636
rect 20772 9596 20778 9608
rect 23106 9596 23112 9608
rect 23164 9596 23170 9648
rect 23750 9636 23756 9648
rect 23711 9608 23756 9636
rect 23750 9596 23756 9608
rect 23808 9596 23814 9648
rect 24118 9596 24124 9648
rect 24176 9636 24182 9648
rect 27890 9636 27896 9648
rect 24176 9608 27896 9636
rect 24176 9596 24182 9608
rect 27890 9596 27896 9608
rect 27948 9596 27954 9648
rect 33229 9639 33287 9645
rect 33229 9605 33241 9639
rect 33275 9636 33287 9639
rect 33502 9636 33508 9648
rect 33275 9608 33508 9636
rect 33275 9605 33287 9608
rect 33229 9599 33287 9605
rect 33502 9596 33508 9608
rect 33560 9596 33566 9648
rect 36262 9596 36268 9648
rect 36320 9636 36326 9648
rect 37016 9636 37044 9667
rect 44358 9664 44364 9716
rect 44416 9713 44422 9716
rect 44416 9707 44465 9713
rect 44416 9673 44419 9707
rect 44453 9673 44465 9707
rect 44416 9667 44465 9673
rect 44545 9707 44603 9713
rect 44545 9673 44557 9707
rect 44591 9704 44603 9707
rect 44910 9704 44916 9716
rect 44591 9676 44916 9704
rect 44591 9673 44603 9676
rect 44545 9667 44603 9673
rect 44416 9664 44422 9667
rect 44910 9664 44916 9676
rect 44968 9704 44974 9716
rect 45186 9704 45192 9716
rect 44968 9676 45192 9704
rect 44968 9664 44974 9676
rect 45186 9664 45192 9676
rect 45244 9664 45250 9716
rect 48130 9664 48136 9716
rect 48188 9704 48194 9716
rect 48590 9704 48596 9716
rect 48188 9676 48596 9704
rect 48188 9664 48194 9676
rect 48590 9664 48596 9676
rect 48648 9664 48654 9716
rect 49050 9704 49056 9716
rect 49011 9676 49056 9704
rect 49050 9664 49056 9676
rect 49108 9664 49114 9716
rect 49988 9676 50936 9704
rect 36320 9608 37044 9636
rect 36320 9596 36326 9608
rect 37090 9596 37096 9648
rect 37148 9636 37154 9648
rect 37148 9608 41828 9636
rect 37148 9596 37154 9608
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9568 18935 9571
rect 19518 9568 19524 9580
rect 18923 9540 19524 9568
rect 18923 9537 18935 9540
rect 18877 9531 18935 9537
rect 19518 9528 19524 9540
rect 19576 9528 19582 9580
rect 22741 9571 22799 9577
rect 19628 9540 22324 9568
rect 18322 9500 18328 9512
rect 16899 9472 17632 9500
rect 18283 9472 18328 9500
rect 16899 9469 16911 9472
rect 16853 9463 16911 9469
rect 18322 9460 18328 9472
rect 18380 9460 18386 9512
rect 18414 9460 18420 9512
rect 18472 9500 18478 9512
rect 19628 9500 19656 9540
rect 18472 9472 19656 9500
rect 18472 9460 18478 9472
rect 19702 9460 19708 9512
rect 19760 9500 19766 9512
rect 19981 9503 20039 9509
rect 19760 9472 19805 9500
rect 19760 9460 19766 9472
rect 19981 9469 19993 9503
rect 20027 9500 20039 9503
rect 20898 9500 20904 9512
rect 20027 9472 20904 9500
rect 20027 9469 20039 9472
rect 19981 9463 20039 9469
rect 20898 9460 20904 9472
rect 20956 9460 20962 9512
rect 21726 9500 21732 9512
rect 21008 9472 21732 9500
rect 21008 9432 21036 9472
rect 21726 9460 21732 9472
rect 21784 9460 21790 9512
rect 22186 9500 22192 9512
rect 22147 9472 22192 9500
rect 22186 9460 22192 9472
rect 22244 9460 22250 9512
rect 22296 9509 22324 9540
rect 22741 9537 22753 9571
rect 22787 9568 22799 9571
rect 23934 9568 23940 9580
rect 22787 9540 23940 9568
rect 22787 9537 22799 9540
rect 22741 9531 22799 9537
rect 23934 9528 23940 9540
rect 23992 9528 23998 9580
rect 26142 9568 26148 9580
rect 25516 9540 26148 9568
rect 22281 9503 22339 9509
rect 22281 9469 22293 9503
rect 22327 9500 22339 9503
rect 23198 9500 23204 9512
rect 22327 9472 23204 9500
rect 22327 9469 22339 9472
rect 22281 9463 22339 9469
rect 23198 9460 23204 9472
rect 23256 9460 23262 9512
rect 23661 9503 23719 9509
rect 23661 9469 23673 9503
rect 23707 9500 23719 9503
rect 24210 9500 24216 9512
rect 23707 9472 24216 9500
rect 23707 9469 23719 9472
rect 23661 9463 23719 9469
rect 24210 9460 24216 9472
rect 24268 9460 24274 9512
rect 25314 9500 25320 9512
rect 25275 9472 25320 9500
rect 25314 9460 25320 9472
rect 25372 9460 25378 9512
rect 25516 9509 25544 9540
rect 26142 9528 26148 9540
rect 26200 9528 26206 9580
rect 26418 9528 26424 9580
rect 26476 9568 26482 9580
rect 26697 9571 26755 9577
rect 26697 9568 26709 9571
rect 26476 9540 26709 9568
rect 26476 9528 26482 9540
rect 26697 9537 26709 9540
rect 26743 9537 26755 9571
rect 26697 9531 26755 9537
rect 27154 9528 27160 9580
rect 27212 9568 27218 9580
rect 29730 9568 29736 9580
rect 27212 9540 29592 9568
rect 29691 9540 29736 9568
rect 27212 9528 27218 9540
rect 25501 9503 25559 9509
rect 25501 9469 25513 9503
rect 25547 9469 25559 9503
rect 25501 9463 25559 9469
rect 25869 9503 25927 9509
rect 25869 9469 25881 9503
rect 25915 9500 25927 9503
rect 27246 9500 27252 9512
rect 25915 9472 27252 9500
rect 25915 9469 25927 9472
rect 25869 9463 25927 9469
rect 27246 9460 27252 9472
rect 27304 9460 27310 9512
rect 27433 9503 27491 9509
rect 27433 9469 27445 9503
rect 27479 9500 27491 9503
rect 27522 9500 27528 9512
rect 27479 9472 27528 9500
rect 27479 9469 27491 9472
rect 27433 9463 27491 9469
rect 27522 9460 27528 9472
rect 27580 9460 27586 9512
rect 27632 9509 27660 9540
rect 27617 9503 27675 9509
rect 27617 9469 27629 9503
rect 27663 9469 27675 9503
rect 27617 9463 27675 9469
rect 27801 9503 27859 9509
rect 27801 9469 27813 9503
rect 27847 9469 27859 9503
rect 27801 9463 27859 9469
rect 28169 9503 28227 9509
rect 28169 9469 28181 9503
rect 28215 9500 28227 9503
rect 28994 9500 29000 9512
rect 28215 9472 29000 9500
rect 28215 9469 28227 9472
rect 28169 9463 28227 9469
rect 14752 9404 19472 9432
rect 8720 9336 9628 9364
rect 8720 9324 8726 9336
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 11333 9367 11391 9373
rect 11333 9364 11345 9367
rect 9732 9336 11345 9364
rect 9732 9324 9738 9336
rect 11333 9333 11345 9336
rect 11379 9364 11391 9367
rect 11790 9364 11796 9376
rect 11379 9336 11796 9364
rect 11379 9333 11391 9336
rect 11333 9327 11391 9333
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 18322 9324 18328 9376
rect 18380 9364 18386 9376
rect 19334 9364 19340 9376
rect 18380 9336 19340 9364
rect 18380 9324 18386 9336
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 19444 9364 19472 9404
rect 20640 9404 21036 9432
rect 20640 9364 20668 9404
rect 21082 9392 21088 9444
rect 21140 9432 21146 9444
rect 21361 9435 21419 9441
rect 21361 9432 21373 9435
rect 21140 9404 21373 9432
rect 21140 9392 21146 9404
rect 21361 9401 21373 9404
rect 21407 9432 21419 9435
rect 22002 9432 22008 9444
rect 21407 9404 22008 9432
rect 21407 9401 21419 9404
rect 21361 9395 21419 9401
rect 22002 9392 22008 9404
rect 22060 9392 22066 9444
rect 26510 9392 26516 9444
rect 26568 9432 26574 9444
rect 27062 9432 27068 9444
rect 26568 9404 27068 9432
rect 26568 9392 26574 9404
rect 27062 9392 27068 9404
rect 27120 9432 27126 9444
rect 27816 9432 27844 9463
rect 28994 9460 29000 9472
rect 29052 9500 29058 9512
rect 29457 9503 29515 9509
rect 29457 9500 29469 9503
rect 29052 9472 29469 9500
rect 29052 9460 29058 9472
rect 29457 9469 29469 9472
rect 29503 9469 29515 9503
rect 29564 9500 29592 9540
rect 29730 9528 29736 9540
rect 29788 9528 29794 9580
rect 32398 9528 32404 9580
rect 32456 9568 32462 9580
rect 37274 9568 37280 9580
rect 32456 9540 37280 9568
rect 32456 9528 32462 9540
rect 37274 9528 37280 9540
rect 37332 9528 37338 9580
rect 39577 9571 39635 9577
rect 39577 9537 39589 9571
rect 39623 9568 39635 9571
rect 41506 9568 41512 9580
rect 39623 9540 41512 9568
rect 39623 9537 39635 9540
rect 39577 9531 39635 9537
rect 41506 9528 41512 9540
rect 41564 9528 41570 9580
rect 41800 9568 41828 9608
rect 42794 9596 42800 9648
rect 42852 9636 42858 9648
rect 48498 9636 48504 9648
rect 42852 9608 48504 9636
rect 42852 9596 42858 9608
rect 48498 9596 48504 9608
rect 48556 9596 48562 9648
rect 48682 9596 48688 9648
rect 48740 9636 48746 9648
rect 49988 9636 50016 9676
rect 48740 9608 50016 9636
rect 50065 9639 50123 9645
rect 48740 9596 48746 9608
rect 50065 9605 50077 9639
rect 50111 9636 50123 9639
rect 50111 9608 50568 9636
rect 50111 9605 50123 9608
rect 50065 9599 50123 9605
rect 43254 9568 43260 9580
rect 41800 9540 43260 9568
rect 43254 9528 43260 9540
rect 43312 9528 43318 9580
rect 43441 9571 43499 9577
rect 43441 9537 43453 9571
rect 43487 9568 43499 9571
rect 43898 9568 43904 9580
rect 43487 9540 43904 9568
rect 43487 9537 43499 9540
rect 43441 9531 43499 9537
rect 43898 9528 43904 9540
rect 43956 9568 43962 9580
rect 44637 9571 44695 9577
rect 44637 9568 44649 9571
rect 43956 9540 44649 9568
rect 43956 9528 43962 9540
rect 44637 9537 44649 9540
rect 44683 9568 44695 9571
rect 45554 9568 45560 9580
rect 44683 9540 45560 9568
rect 44683 9537 44695 9540
rect 44637 9531 44695 9537
rect 45554 9528 45560 9540
rect 45612 9528 45618 9580
rect 46106 9568 46112 9580
rect 46067 9540 46112 9568
rect 46106 9528 46112 9540
rect 46164 9528 46170 9580
rect 48225 9571 48283 9577
rect 48225 9568 48237 9571
rect 46216 9540 48237 9568
rect 29564 9472 31800 9500
rect 29457 9463 29515 9469
rect 29270 9432 29276 9444
rect 27120 9404 27844 9432
rect 29231 9404 29276 9432
rect 27120 9392 27126 9404
rect 29270 9392 29276 9404
rect 29328 9392 29334 9444
rect 30742 9432 30748 9444
rect 30703 9404 30748 9432
rect 30742 9392 30748 9404
rect 30800 9392 30806 9444
rect 31772 9432 31800 9472
rect 31846 9460 31852 9512
rect 31904 9500 31910 9512
rect 32585 9503 32643 9509
rect 32585 9500 32597 9503
rect 31904 9472 32597 9500
rect 31904 9460 31910 9472
rect 32585 9469 32597 9472
rect 32631 9500 32643 9503
rect 32674 9500 32680 9512
rect 32631 9472 32680 9500
rect 32631 9469 32643 9472
rect 32585 9463 32643 9469
rect 32674 9460 32680 9472
rect 32732 9460 32738 9512
rect 33410 9500 33416 9512
rect 33371 9472 33416 9500
rect 33410 9460 33416 9472
rect 33468 9460 33474 9512
rect 33781 9503 33839 9509
rect 33781 9469 33793 9503
rect 33827 9469 33839 9503
rect 33781 9463 33839 9469
rect 33796 9432 33824 9463
rect 33870 9460 33876 9512
rect 33928 9500 33934 9512
rect 35342 9500 35348 9512
rect 33928 9472 35112 9500
rect 35303 9472 35348 9500
rect 33928 9460 33934 9472
rect 33962 9432 33968 9444
rect 31772 9404 33732 9432
rect 33796 9404 33968 9432
rect 19444 9336 20668 9364
rect 20990 9324 20996 9376
rect 21048 9364 21054 9376
rect 21634 9364 21640 9376
rect 21048 9336 21640 9364
rect 21048 9324 21054 9336
rect 21634 9324 21640 9336
rect 21692 9364 21698 9376
rect 27798 9364 27804 9376
rect 21692 9336 27804 9364
rect 21692 9324 21698 9336
rect 27798 9324 27804 9336
rect 27856 9324 27862 9376
rect 31294 9324 31300 9376
rect 31352 9364 31358 9376
rect 32033 9367 32091 9373
rect 32033 9364 32045 9367
rect 31352 9336 32045 9364
rect 31352 9324 31358 9336
rect 32033 9333 32045 9336
rect 32079 9364 32091 9367
rect 32398 9364 32404 9376
rect 32079 9336 32404 9364
rect 32079 9333 32091 9336
rect 32033 9327 32091 9333
rect 32398 9324 32404 9336
rect 32456 9324 32462 9376
rect 32766 9364 32772 9376
rect 32727 9336 32772 9364
rect 32766 9324 32772 9336
rect 32824 9324 32830 9376
rect 33704 9364 33732 9404
rect 33962 9392 33968 9404
rect 34020 9392 34026 9444
rect 34885 9435 34943 9441
rect 34885 9401 34897 9435
rect 34931 9432 34943 9435
rect 34974 9432 34980 9444
rect 34931 9404 34980 9432
rect 34931 9401 34943 9404
rect 34885 9395 34943 9401
rect 34974 9392 34980 9404
rect 35032 9392 35038 9444
rect 34790 9364 34796 9376
rect 33704 9336 34796 9364
rect 34790 9324 34796 9336
rect 34848 9324 34854 9376
rect 35084 9364 35112 9472
rect 35342 9460 35348 9472
rect 35400 9460 35406 9512
rect 35434 9460 35440 9512
rect 35492 9500 35498 9512
rect 35529 9503 35587 9509
rect 35529 9500 35541 9503
rect 35492 9472 35541 9500
rect 35492 9460 35498 9472
rect 35529 9469 35541 9472
rect 35575 9469 35587 9503
rect 35529 9463 35587 9469
rect 35713 9503 35771 9509
rect 35713 9469 35725 9503
rect 35759 9500 35771 9503
rect 35894 9500 35900 9512
rect 35759 9472 35900 9500
rect 35759 9469 35771 9472
rect 35713 9463 35771 9469
rect 35894 9460 35900 9472
rect 35952 9460 35958 9512
rect 36446 9460 36452 9512
rect 36504 9500 36510 9512
rect 36722 9500 36728 9512
rect 36504 9472 36728 9500
rect 36504 9460 36510 9472
rect 36722 9460 36728 9472
rect 36780 9460 36786 9512
rect 36817 9503 36875 9509
rect 36817 9469 36829 9503
rect 36863 9469 36875 9503
rect 36817 9463 36875 9469
rect 36630 9392 36636 9444
rect 36688 9432 36694 9444
rect 36832 9432 36860 9463
rect 38746 9460 38752 9512
rect 38804 9500 38810 9512
rect 39025 9503 39083 9509
rect 39025 9500 39037 9503
rect 38804 9472 39037 9500
rect 38804 9460 38810 9472
rect 39025 9469 39037 9472
rect 39071 9469 39083 9503
rect 39025 9463 39083 9469
rect 39117 9503 39175 9509
rect 39117 9469 39129 9503
rect 39163 9469 39175 9503
rect 41414 9500 41420 9512
rect 41375 9472 41420 9500
rect 39117 9463 39175 9469
rect 37274 9432 37280 9444
rect 36688 9404 37280 9432
rect 36688 9392 36694 9404
rect 37274 9392 37280 9404
rect 37332 9392 37338 9444
rect 36814 9364 36820 9376
rect 35084 9336 36820 9364
rect 36814 9324 36820 9336
rect 36872 9324 36878 9376
rect 39040 9364 39068 9463
rect 39132 9432 39160 9463
rect 41414 9460 41420 9472
rect 41472 9460 41478 9512
rect 41785 9503 41843 9509
rect 41785 9469 41797 9503
rect 41831 9500 41843 9503
rect 41874 9500 41880 9512
rect 41831 9472 41880 9500
rect 41831 9469 41843 9472
rect 41785 9463 41843 9469
rect 41874 9460 41880 9472
rect 41932 9460 41938 9512
rect 42058 9500 42064 9512
rect 42019 9472 42064 9500
rect 42058 9460 42064 9472
rect 42116 9460 42122 9512
rect 44358 9460 44364 9512
rect 44416 9500 44422 9512
rect 46216 9500 46244 9540
rect 48225 9537 48237 9540
rect 48271 9537 48283 9571
rect 48225 9531 48283 9537
rect 46382 9500 46388 9512
rect 44416 9472 46244 9500
rect 46343 9472 46388 9500
rect 44416 9460 44422 9472
rect 46382 9460 46388 9472
rect 46440 9460 46446 9512
rect 47486 9460 47492 9512
rect 47544 9500 47550 9512
rect 47673 9503 47731 9509
rect 47673 9500 47685 9503
rect 47544 9472 47685 9500
rect 47544 9460 47550 9472
rect 47673 9469 47685 9472
rect 47719 9469 47731 9503
rect 47673 9463 47731 9469
rect 47762 9460 47768 9512
rect 47820 9500 47826 9512
rect 49234 9500 49240 9512
rect 47820 9472 47865 9500
rect 49195 9472 49240 9500
rect 47820 9460 47826 9472
rect 49234 9460 49240 9472
rect 49292 9460 49298 9512
rect 49786 9460 49792 9512
rect 49844 9500 49850 9512
rect 50249 9503 50307 9509
rect 50249 9500 50261 9503
rect 49844 9472 50261 9500
rect 49844 9460 49850 9472
rect 50249 9469 50261 9472
rect 50295 9469 50307 9503
rect 50430 9500 50436 9512
rect 50391 9472 50436 9500
rect 50249 9463 50307 9469
rect 50430 9460 50436 9472
rect 50488 9460 50494 9512
rect 39298 9432 39304 9444
rect 39132 9404 39304 9432
rect 39298 9392 39304 9404
rect 39356 9392 39362 9444
rect 44082 9432 44088 9444
rect 43272 9404 44088 9432
rect 39942 9364 39948 9376
rect 39040 9336 39948 9364
rect 39942 9324 39948 9336
rect 40000 9324 40006 9376
rect 41233 9367 41291 9373
rect 41233 9333 41245 9367
rect 41279 9364 41291 9367
rect 43272 9364 43300 9404
rect 44082 9392 44088 9404
rect 44140 9392 44146 9444
rect 44269 9435 44327 9441
rect 44269 9401 44281 9435
rect 44315 9432 44327 9435
rect 46106 9432 46112 9444
rect 44315 9404 46112 9432
rect 44315 9401 44327 9404
rect 44269 9395 44327 9401
rect 46106 9392 46112 9404
rect 46164 9392 46170 9444
rect 46474 9392 46480 9444
rect 46532 9432 46538 9444
rect 46842 9432 46848 9444
rect 46532 9404 46625 9432
rect 46803 9404 46848 9432
rect 46532 9392 46538 9404
rect 46842 9392 46848 9404
rect 46900 9392 46906 9444
rect 50540 9432 50568 9608
rect 50908 9568 50936 9676
rect 54846 9636 54852 9648
rect 54588 9608 54852 9636
rect 54588 9568 54616 9608
rect 54846 9596 54852 9608
rect 54904 9596 54910 9648
rect 50908 9540 54616 9568
rect 54662 9528 54668 9580
rect 54720 9568 54726 9580
rect 59449 9571 59507 9577
rect 59449 9568 59461 9571
rect 54720 9540 59461 9568
rect 54720 9528 54726 9540
rect 59449 9537 59461 9540
rect 59495 9537 59507 9571
rect 59449 9531 59507 9537
rect 50617 9503 50675 9509
rect 50617 9469 50629 9503
rect 50663 9500 50675 9503
rect 51258 9500 51264 9512
rect 50663 9472 51264 9500
rect 50663 9469 50675 9472
rect 50617 9463 50675 9469
rect 51258 9460 51264 9472
rect 51316 9460 51322 9512
rect 51534 9460 51540 9512
rect 51592 9500 51598 9512
rect 52641 9503 52699 9509
rect 52641 9500 52653 9503
rect 51592 9472 52653 9500
rect 51592 9460 51598 9472
rect 52641 9469 52653 9472
rect 52687 9469 52699 9503
rect 52641 9463 52699 9469
rect 52730 9460 52736 9512
rect 52788 9500 52794 9512
rect 52917 9503 52975 9509
rect 52917 9500 52929 9503
rect 52788 9472 52929 9500
rect 52788 9460 52794 9472
rect 52917 9469 52929 9472
rect 52963 9469 52975 9503
rect 52917 9463 52975 9469
rect 54846 9460 54852 9512
rect 54904 9500 54910 9512
rect 55401 9503 55459 9509
rect 55401 9500 55413 9503
rect 54904 9472 55413 9500
rect 54904 9460 54910 9472
rect 55401 9469 55413 9472
rect 55447 9469 55459 9503
rect 55401 9463 55459 9469
rect 51718 9432 51724 9444
rect 50540 9404 51724 9432
rect 51718 9392 51724 9404
rect 51776 9392 51782 9444
rect 54754 9392 54760 9444
rect 54812 9432 54818 9444
rect 55217 9435 55275 9441
rect 55217 9432 55229 9435
rect 54812 9404 55229 9432
rect 54812 9392 54818 9404
rect 55217 9401 55229 9404
rect 55263 9401 55275 9435
rect 55217 9395 55275 9401
rect 41279 9336 43300 9364
rect 41279 9333 41291 9336
rect 41233 9327 41291 9333
rect 43346 9324 43352 9376
rect 43404 9364 43410 9376
rect 44913 9367 44971 9373
rect 44913 9364 44925 9367
rect 43404 9336 44925 9364
rect 43404 9324 43410 9336
rect 44913 9333 44925 9336
rect 44959 9333 44971 9367
rect 44913 9327 44971 9333
rect 45002 9324 45008 9376
rect 45060 9364 45066 9376
rect 46198 9364 46204 9376
rect 45060 9336 46204 9364
rect 45060 9324 45066 9336
rect 46198 9324 46204 9336
rect 46256 9364 46262 9376
rect 46293 9367 46351 9373
rect 46293 9364 46305 9367
rect 46256 9336 46305 9364
rect 46256 9324 46262 9336
rect 46293 9333 46305 9336
rect 46339 9333 46351 9367
rect 46492 9364 46520 9392
rect 49418 9364 49424 9376
rect 46492 9336 49424 9364
rect 46293 9327 46351 9333
rect 49418 9324 49424 9336
rect 49476 9324 49482 9376
rect 52914 9324 52920 9376
rect 52972 9364 52978 9376
rect 54021 9367 54079 9373
rect 54021 9364 54033 9367
rect 52972 9336 54033 9364
rect 52972 9324 52978 9336
rect 54021 9333 54033 9336
rect 54067 9364 54079 9367
rect 54294 9364 54300 9376
rect 54067 9336 54300 9364
rect 54067 9333 54079 9336
rect 54021 9327 54079 9333
rect 54294 9324 54300 9336
rect 54352 9324 54358 9376
rect 55416 9364 55444 9463
rect 57330 9460 57336 9512
rect 57388 9500 57394 9512
rect 57974 9500 57980 9512
rect 57388 9472 57980 9500
rect 57388 9460 57394 9472
rect 57974 9460 57980 9472
rect 58032 9500 58038 9512
rect 58069 9503 58127 9509
rect 58069 9500 58081 9503
rect 58032 9472 58081 9500
rect 58032 9460 58038 9472
rect 58069 9469 58081 9472
rect 58115 9469 58127 9503
rect 58342 9500 58348 9512
rect 58303 9472 58348 9500
rect 58069 9463 58127 9469
rect 58342 9460 58348 9472
rect 58400 9460 58406 9512
rect 55766 9432 55772 9444
rect 55727 9404 55772 9432
rect 55766 9392 55772 9404
rect 55824 9392 55830 9444
rect 60182 9364 60188 9376
rect 55416 9336 60188 9364
rect 60182 9324 60188 9336
rect 60240 9324 60246 9376
rect 1104 9274 62192 9296
rect 1104 9222 21344 9274
rect 21396 9222 21408 9274
rect 21460 9222 21472 9274
rect 21524 9222 21536 9274
rect 21588 9222 41707 9274
rect 41759 9222 41771 9274
rect 41823 9222 41835 9274
rect 41887 9222 41899 9274
rect 41951 9222 62192 9274
rect 1104 9200 62192 9222
rect 382 9120 388 9172
rect 440 9160 446 9172
rect 30742 9160 30748 9172
rect 440 9132 30748 9160
rect 440 9120 446 9132
rect 30742 9120 30748 9132
rect 30800 9120 30806 9172
rect 32306 9120 32312 9172
rect 32364 9160 32370 9172
rect 36630 9160 36636 9172
rect 32364 9132 36636 9160
rect 32364 9120 32370 9132
rect 36630 9120 36636 9132
rect 36688 9120 36694 9172
rect 36722 9120 36728 9172
rect 36780 9160 36786 9172
rect 58342 9160 58348 9172
rect 36780 9132 51948 9160
rect 36780 9120 36786 9132
rect 2133 9095 2191 9101
rect 2133 9061 2145 9095
rect 2179 9092 2191 9095
rect 3234 9092 3240 9104
rect 2179 9064 3240 9092
rect 2179 9061 2191 9064
rect 2133 9055 2191 9061
rect 3234 9052 3240 9064
rect 3292 9052 3298 9104
rect 4706 9092 4712 9104
rect 4667 9064 4712 9092
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 9582 9092 9588 9104
rect 8220 9064 9588 9092
rect 2593 9027 2651 9033
rect 2593 8993 2605 9027
rect 2639 9024 2651 9027
rect 2866 9024 2872 9036
rect 2639 8996 2872 9024
rect 2639 8993 2651 8996
rect 2593 8987 2651 8993
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 2958 8984 2964 9036
rect 3016 9024 3022 9036
rect 3016 8996 3061 9024
rect 3016 8984 3022 8996
rect 4522 8984 4528 9036
rect 4580 9024 4586 9036
rect 5169 9027 5227 9033
rect 5169 9024 5181 9027
rect 4580 8996 5181 9024
rect 4580 8984 4586 8996
rect 5169 8993 5181 8996
rect 5215 8993 5227 9027
rect 5534 9024 5540 9036
rect 5495 8996 5540 9024
rect 5169 8987 5227 8993
rect 5534 8984 5540 8996
rect 5592 8984 5598 9036
rect 5626 8984 5632 9036
rect 5684 9024 5690 9036
rect 7466 9024 7472 9036
rect 5684 8996 7472 9024
rect 5684 8984 5690 8996
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 8220 8968 8248 9064
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 10336 9064 10824 9092
rect 10336 9033 10364 9064
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 8993 8355 9027
rect 8297 8987 8355 8993
rect 10321 9027 10379 9033
rect 10321 8993 10333 9027
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 3050 8956 3056 8968
rect 3011 8928 3056 8956
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 8202 8956 8208 8968
rect 8163 8928 8208 8956
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 8312 8888 8340 8987
rect 10594 8984 10600 9036
rect 10652 9024 10658 9036
rect 10689 9027 10747 9033
rect 10689 9024 10701 9027
rect 10652 8996 10701 9024
rect 10652 8984 10658 8996
rect 10689 8993 10701 8996
rect 10735 8993 10747 9027
rect 10796 9024 10824 9064
rect 11790 9052 11796 9104
rect 11848 9092 11854 9104
rect 14274 9092 14280 9104
rect 11848 9064 12756 9092
rect 11848 9052 11854 9064
rect 12342 9024 12348 9036
rect 10796 8996 12348 9024
rect 10689 8987 10747 8993
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 12728 9033 12756 9064
rect 12912 9064 14280 9092
rect 12912 9033 12940 9064
rect 12713 9027 12771 9033
rect 12713 8993 12725 9027
rect 12759 8993 12771 9027
rect 12713 8987 12771 8993
rect 12897 9027 12955 9033
rect 12897 8993 12909 9027
rect 12943 8993 12955 9027
rect 13722 9024 13728 9036
rect 13683 8996 13728 9024
rect 12897 8987 12955 8993
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 8803 8928 10241 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 10778 8956 10784 8968
rect 10739 8928 10784 8956
rect 10229 8919 10287 8925
rect 10778 8916 10784 8928
rect 10836 8916 10842 8968
rect 11054 8916 11060 8968
rect 11112 8956 11118 8968
rect 11701 8959 11759 8965
rect 11701 8956 11713 8959
rect 11112 8928 11713 8956
rect 11112 8916 11118 8928
rect 11701 8925 11713 8928
rect 11747 8925 11759 8959
rect 12250 8956 12256 8968
rect 12211 8928 12256 8956
rect 11701 8919 11759 8925
rect 12250 8916 12256 8928
rect 12308 8916 12314 8968
rect 8312 8860 9904 8888
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 9769 8823 9827 8829
rect 9769 8820 9781 8823
rect 8444 8792 9781 8820
rect 8444 8780 8450 8792
rect 9769 8789 9781 8792
rect 9815 8789 9827 8823
rect 9876 8820 9904 8860
rect 12912 8820 12940 8987
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 13924 9033 13952 9064
rect 14274 9052 14280 9064
rect 14332 9092 14338 9104
rect 17034 9092 17040 9104
rect 14332 9064 16712 9092
rect 16995 9064 17040 9092
rect 14332 9052 14338 9064
rect 13909 9027 13967 9033
rect 13909 8993 13921 9027
rect 13955 8993 13967 9027
rect 13909 8987 13967 8993
rect 16209 9027 16267 9033
rect 16209 8993 16221 9027
rect 16255 9024 16267 9027
rect 16390 9024 16396 9036
rect 16255 8996 16396 9024
rect 16255 8993 16267 8996
rect 16209 8987 16267 8993
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 16577 9027 16635 9033
rect 16577 8993 16589 9027
rect 16623 8993 16635 9027
rect 16684 9024 16712 9064
rect 17034 9052 17040 9064
rect 17092 9052 17098 9104
rect 18690 9052 18696 9104
rect 18748 9092 18754 9104
rect 20714 9092 20720 9104
rect 18748 9064 20720 9092
rect 18748 9052 18754 9064
rect 17957 9027 18015 9033
rect 17957 9024 17969 9027
rect 16684 8996 17969 9024
rect 16577 8987 16635 8993
rect 17957 8993 17969 8996
rect 18003 8993 18015 9027
rect 17957 8987 18015 8993
rect 16482 8956 16488 8968
rect 16443 8928 16488 8956
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 16592 8956 16620 8987
rect 18506 8984 18512 9036
rect 18564 9024 18570 9036
rect 19444 9033 19472 9064
rect 20714 9052 20720 9064
rect 20772 9052 20778 9104
rect 20898 9092 20904 9104
rect 20859 9064 20904 9092
rect 20898 9052 20904 9064
rect 20956 9052 20962 9104
rect 21818 9052 21824 9104
rect 21876 9092 21882 9104
rect 23293 9095 23351 9101
rect 23293 9092 23305 9095
rect 21876 9064 23305 9092
rect 21876 9052 21882 9064
rect 23293 9061 23305 9064
rect 23339 9061 23351 9095
rect 23293 9055 23351 9061
rect 24857 9095 24915 9101
rect 24857 9061 24869 9095
rect 24903 9092 24915 9095
rect 24946 9092 24952 9104
rect 24903 9064 24952 9092
rect 24903 9061 24915 9064
rect 24857 9055 24915 9061
rect 24946 9052 24952 9064
rect 25004 9052 25010 9104
rect 28721 9095 28779 9101
rect 28721 9061 28733 9095
rect 28767 9092 28779 9095
rect 28902 9092 28908 9104
rect 28767 9064 28908 9092
rect 28767 9061 28779 9064
rect 28721 9055 28779 9061
rect 19245 9027 19303 9033
rect 19245 9024 19257 9027
rect 18564 8996 19257 9024
rect 18564 8984 18570 8996
rect 19245 8993 19257 8996
rect 19291 8993 19303 9027
rect 19245 8987 19303 8993
rect 19392 9027 19472 9033
rect 19392 8993 19404 9027
rect 19438 8996 19472 9027
rect 19536 8996 21496 9024
rect 19438 8993 19450 8996
rect 19392 8987 19450 8993
rect 17770 8956 17776 8968
rect 16592 8928 17776 8956
rect 9876 8792 12940 8820
rect 9769 8783 9827 8789
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 14001 8823 14059 8829
rect 14001 8820 14013 8823
rect 13872 8792 14013 8820
rect 13872 8780 13878 8792
rect 14001 8789 14013 8792
rect 14047 8789 14059 8823
rect 14001 8783 14059 8789
rect 15930 8780 15936 8832
rect 15988 8820 15994 8832
rect 16025 8823 16083 8829
rect 16025 8820 16037 8823
rect 15988 8792 16037 8820
rect 15988 8780 15994 8792
rect 16025 8789 16037 8792
rect 16071 8789 16083 8823
rect 16025 8783 16083 8789
rect 16114 8780 16120 8832
rect 16172 8820 16178 8832
rect 16684 8820 16712 8928
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8925 17923 8959
rect 17865 8919 17923 8925
rect 18417 8959 18475 8965
rect 18417 8925 18429 8959
rect 18463 8956 18475 8959
rect 19536 8956 19564 8996
rect 18463 8928 19564 8956
rect 18463 8925 18475 8928
rect 18417 8919 18475 8925
rect 16172 8792 16712 8820
rect 17880 8820 17908 8919
rect 19610 8916 19616 8968
rect 19668 8956 19674 8968
rect 19668 8928 19713 8956
rect 19668 8916 19674 8928
rect 20070 8916 20076 8968
rect 20128 8956 20134 8968
rect 21174 8956 21180 8968
rect 20128 8928 21180 8956
rect 20128 8916 20134 8928
rect 21174 8916 21180 8928
rect 21232 8916 21238 8968
rect 21468 8965 21496 8996
rect 21542 8984 21548 9036
rect 21600 9024 21606 9036
rect 21913 9027 21971 9033
rect 21600 8996 21645 9024
rect 21600 8984 21606 8996
rect 21913 8993 21925 9027
rect 21959 9024 21971 9027
rect 22278 9024 22284 9036
rect 21959 8996 22284 9024
rect 21959 8993 21971 8996
rect 21913 8987 21971 8993
rect 22278 8984 22284 8996
rect 22336 8984 22342 9036
rect 23106 9024 23112 9036
rect 23067 8996 23112 9024
rect 23106 8984 23112 8996
rect 23164 8984 23170 9036
rect 23201 9027 23259 9033
rect 23201 8993 23213 9027
rect 23247 8993 23259 9027
rect 24762 9024 24768 9036
rect 24723 8996 24768 9024
rect 23201 8987 23259 8993
rect 21453 8959 21511 8965
rect 21453 8925 21465 8959
rect 21499 8925 21511 8959
rect 21453 8919 21511 8925
rect 21818 8916 21824 8968
rect 21876 8956 21882 8968
rect 22005 8959 22063 8965
rect 22005 8956 22017 8959
rect 21876 8928 22017 8956
rect 21876 8916 21882 8928
rect 22005 8925 22017 8928
rect 22051 8925 22063 8959
rect 22005 8919 22063 8925
rect 22094 8916 22100 8968
rect 22152 8956 22158 8968
rect 22925 8959 22983 8965
rect 22925 8956 22937 8959
rect 22152 8928 22937 8956
rect 22152 8916 22158 8928
rect 22925 8925 22937 8928
rect 22971 8925 22983 8959
rect 23216 8956 23244 8987
rect 24762 8984 24768 8996
rect 24820 8984 24826 9036
rect 27798 8984 27804 9036
rect 27856 9024 27862 9036
rect 28736 9024 28764 9055
rect 28902 9052 28908 9064
rect 28960 9052 28966 9104
rect 35618 9092 35624 9104
rect 35579 9064 35624 9092
rect 35618 9052 35624 9064
rect 35676 9052 35682 9104
rect 37090 9092 37096 9104
rect 35912 9064 37096 9092
rect 27856 8996 28764 9024
rect 27856 8984 27862 8996
rect 29178 8984 29184 9036
rect 29236 9024 29242 9036
rect 30009 9027 30067 9033
rect 30009 9024 30021 9027
rect 29236 8996 30021 9024
rect 29236 8984 29242 8996
rect 30009 8993 30021 8996
rect 30055 8993 30067 9027
rect 30650 9024 30656 9036
rect 30611 8996 30656 9024
rect 30009 8987 30067 8993
rect 30650 8984 30656 8996
rect 30708 8984 30714 9036
rect 32122 9024 32128 9036
rect 32035 8996 32128 9024
rect 32122 8984 32128 8996
rect 32180 9024 32186 9036
rect 32490 9024 32496 9036
rect 32180 8996 32496 9024
rect 32180 8984 32186 8996
rect 32490 8984 32496 8996
rect 32548 8984 32554 9036
rect 34793 9027 34851 9033
rect 34793 8993 34805 9027
rect 34839 9024 34851 9027
rect 34882 9024 34888 9036
rect 34839 8996 34888 9024
rect 34839 8993 34851 8996
rect 34793 8987 34851 8993
rect 34882 8984 34888 8996
rect 34940 9024 34946 9036
rect 35912 9024 35940 9064
rect 37090 9052 37096 9064
rect 37148 9052 37154 9104
rect 38289 9095 38347 9101
rect 38289 9061 38301 9095
rect 38335 9092 38347 9095
rect 38654 9092 38660 9104
rect 38335 9064 38660 9092
rect 38335 9061 38347 9064
rect 38289 9055 38347 9061
rect 38654 9052 38660 9064
rect 38712 9052 38718 9104
rect 39316 9064 40172 9092
rect 39316 9036 39344 9064
rect 36078 9024 36084 9036
rect 34940 8996 35940 9024
rect 36039 8996 36084 9024
rect 34940 8984 34946 8996
rect 36078 8984 36084 8996
rect 36136 8984 36142 9036
rect 36449 9027 36507 9033
rect 36449 8993 36461 9027
rect 36495 8993 36507 9027
rect 36449 8987 36507 8993
rect 36541 9027 36599 9033
rect 36541 8993 36553 9027
rect 36587 9024 36599 9027
rect 36814 9024 36820 9036
rect 36587 8996 36820 9024
rect 36587 8993 36599 8996
rect 36541 8987 36599 8993
rect 23658 8956 23664 8968
rect 22925 8919 22983 8925
rect 23124 8928 23244 8956
rect 23619 8928 23664 8956
rect 17954 8848 17960 8900
rect 18012 8888 18018 8900
rect 22370 8888 22376 8900
rect 18012 8860 22376 8888
rect 18012 8848 18018 8860
rect 22370 8848 22376 8860
rect 22428 8848 22434 8900
rect 22554 8848 22560 8900
rect 22612 8888 22618 8900
rect 22738 8888 22744 8900
rect 22612 8860 22744 8888
rect 22612 8848 22618 8860
rect 22738 8848 22744 8860
rect 22796 8888 22802 8900
rect 23124 8888 23152 8928
rect 23658 8916 23664 8928
rect 23716 8916 23722 8968
rect 24946 8916 24952 8968
rect 25004 8956 25010 8968
rect 27065 8959 27123 8965
rect 27065 8956 27077 8959
rect 25004 8928 27077 8956
rect 25004 8916 25010 8928
rect 27065 8925 27077 8928
rect 27111 8925 27123 8959
rect 27338 8956 27344 8968
rect 27299 8928 27344 8956
rect 27065 8919 27123 8925
rect 27338 8916 27344 8928
rect 27396 8916 27402 8968
rect 27430 8916 27436 8968
rect 27488 8956 27494 8968
rect 31294 8956 31300 8968
rect 27488 8928 31300 8956
rect 27488 8916 27494 8928
rect 31294 8916 31300 8928
rect 31352 8956 31358 8968
rect 32217 8959 32275 8965
rect 32217 8956 32229 8959
rect 31352 8928 32229 8956
rect 31352 8916 31358 8928
rect 32217 8925 32229 8928
rect 32263 8925 32275 8959
rect 32217 8919 32275 8925
rect 32950 8916 32956 8968
rect 33008 8956 33014 8968
rect 33137 8959 33195 8965
rect 33137 8956 33149 8959
rect 33008 8928 33149 8956
rect 33008 8916 33014 8928
rect 33137 8925 33149 8928
rect 33183 8925 33195 8959
rect 33410 8956 33416 8968
rect 33371 8928 33416 8956
rect 33137 8919 33195 8925
rect 33410 8916 33416 8928
rect 33468 8916 33474 8968
rect 35066 8916 35072 8968
rect 35124 8956 35130 8968
rect 36464 8956 36492 8987
rect 36814 8984 36820 8996
rect 36872 8984 36878 9036
rect 37829 9027 37887 9033
rect 37829 8993 37841 9027
rect 37875 9024 37887 9027
rect 39298 9024 39304 9036
rect 37875 8996 39304 9024
rect 37875 8993 37887 8996
rect 37829 8987 37887 8993
rect 39298 8984 39304 8996
rect 39356 8984 39362 9036
rect 39853 9027 39911 9033
rect 39853 8993 39865 9027
rect 39899 8993 39911 9027
rect 39853 8987 39911 8993
rect 35124 8928 36492 8956
rect 35124 8916 35130 8928
rect 36722 8916 36728 8968
rect 36780 8956 36786 8968
rect 37737 8959 37795 8965
rect 37737 8956 37749 8959
rect 36780 8928 37749 8956
rect 36780 8916 36786 8928
rect 37737 8925 37749 8928
rect 37783 8925 37795 8959
rect 37737 8919 37795 8925
rect 22796 8860 23152 8888
rect 22796 8848 22802 8860
rect 23198 8848 23204 8900
rect 23256 8888 23262 8900
rect 23842 8888 23848 8900
rect 23256 8860 23848 8888
rect 23256 8848 23262 8860
rect 23842 8848 23848 8860
rect 23900 8888 23906 8900
rect 36998 8888 37004 8900
rect 23900 8860 26740 8888
rect 23900 8848 23906 8860
rect 19521 8823 19579 8829
rect 19521 8820 19533 8823
rect 17880 8792 19533 8820
rect 16172 8780 16178 8792
rect 19521 8789 19533 8792
rect 19567 8820 19579 8823
rect 19794 8820 19800 8832
rect 19567 8792 19800 8820
rect 19567 8789 19579 8792
rect 19521 8783 19579 8789
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 19889 8823 19947 8829
rect 19889 8789 19901 8823
rect 19935 8820 19947 8823
rect 20806 8820 20812 8832
rect 19935 8792 20812 8820
rect 19935 8789 19947 8792
rect 19889 8783 19947 8789
rect 20806 8780 20812 8792
rect 20864 8780 20870 8832
rect 20898 8780 20904 8832
rect 20956 8820 20962 8832
rect 23382 8820 23388 8832
rect 20956 8792 23388 8820
rect 20956 8780 20962 8792
rect 23382 8780 23388 8792
rect 23440 8780 23446 8832
rect 25406 8780 25412 8832
rect 25464 8820 25470 8832
rect 26602 8820 26608 8832
rect 25464 8792 26608 8820
rect 25464 8780 25470 8792
rect 26602 8780 26608 8792
rect 26660 8780 26666 8832
rect 26712 8820 26740 8860
rect 34072 8860 37004 8888
rect 29730 8820 29736 8832
rect 26712 8792 29736 8820
rect 29730 8780 29736 8792
rect 29788 8780 29794 8832
rect 30190 8820 30196 8832
rect 30151 8792 30196 8820
rect 30190 8780 30196 8792
rect 30248 8780 30254 8832
rect 30558 8780 30564 8832
rect 30616 8820 30622 8832
rect 30837 8823 30895 8829
rect 30837 8820 30849 8823
rect 30616 8792 30849 8820
rect 30616 8780 30622 8792
rect 30837 8789 30849 8792
rect 30883 8789 30895 8823
rect 30837 8783 30895 8789
rect 33042 8780 33048 8832
rect 33100 8820 33106 8832
rect 34072 8820 34100 8860
rect 36998 8848 37004 8860
rect 37056 8848 37062 8900
rect 37918 8888 37924 8900
rect 37108 8860 37924 8888
rect 33100 8792 34100 8820
rect 33100 8780 33106 8792
rect 34790 8780 34796 8832
rect 34848 8820 34854 8832
rect 37108 8820 37136 8860
rect 37918 8848 37924 8860
rect 37976 8888 37982 8900
rect 39868 8888 39896 8987
rect 39942 8984 39948 9036
rect 40000 9024 40006 9036
rect 40037 9027 40095 9033
rect 40037 9024 40049 9027
rect 40000 8996 40049 9024
rect 40000 8984 40006 8996
rect 40037 8993 40049 8996
rect 40083 8993 40095 9027
rect 40144 9024 40172 9064
rect 41598 9052 41604 9104
rect 41656 9092 41662 9104
rect 41785 9095 41843 9101
rect 41785 9092 41797 9095
rect 41656 9064 41797 9092
rect 41656 9052 41662 9064
rect 41785 9061 41797 9064
rect 41831 9061 41843 9095
rect 41785 9055 41843 9061
rect 43254 9052 43260 9104
rect 43312 9092 43318 9104
rect 43312 9064 45048 9092
rect 43312 9052 43318 9064
rect 41325 9027 41383 9033
rect 41325 9024 41337 9027
rect 40144 8996 41337 9024
rect 40037 8987 40095 8993
rect 41325 8993 41337 8996
rect 41371 8993 41383 9027
rect 41325 8987 41383 8993
rect 44177 9027 44235 9033
rect 44177 8993 44189 9027
rect 44223 8993 44235 9027
rect 44177 8987 44235 8993
rect 41233 8959 41291 8965
rect 41233 8925 41245 8959
rect 41279 8925 41291 8959
rect 43990 8956 43996 8968
rect 43951 8928 43996 8956
rect 41233 8919 41291 8925
rect 37976 8860 39896 8888
rect 41248 8888 41276 8919
rect 43990 8916 43996 8928
rect 44048 8916 44054 8968
rect 44192 8956 44220 8987
rect 44266 8984 44272 9036
rect 44324 9024 44330 9036
rect 44729 9027 44787 9033
rect 44729 9024 44741 9027
rect 44324 8996 44741 9024
rect 44324 8984 44330 8996
rect 44729 8993 44741 8996
rect 44775 8993 44787 9027
rect 44910 9024 44916 9036
rect 44871 8996 44916 9024
rect 44729 8987 44787 8993
rect 44910 8984 44916 8996
rect 44968 8984 44974 9036
rect 45020 9024 45048 9064
rect 45646 9052 45652 9104
rect 45704 9092 45710 9104
rect 46385 9095 46443 9101
rect 46385 9092 46397 9095
rect 45704 9064 46397 9092
rect 45704 9052 45710 9064
rect 46385 9061 46397 9064
rect 46431 9061 46443 9095
rect 46385 9055 46443 9061
rect 46569 9095 46627 9101
rect 46569 9061 46581 9095
rect 46615 9092 46627 9095
rect 49421 9095 49479 9101
rect 46615 9064 48820 9092
rect 46615 9061 46627 9064
rect 46569 9055 46627 9061
rect 45020 8996 45140 9024
rect 45112 8956 45140 8996
rect 45462 8984 45468 9036
rect 45520 9024 45526 9036
rect 46477 9027 46535 9033
rect 46477 9024 46489 9027
rect 45520 8996 46489 9024
rect 45520 8984 45526 8996
rect 46477 8993 46489 8996
rect 46523 9024 46535 9027
rect 46523 8996 47900 9024
rect 46523 8993 46535 8996
rect 46477 8987 46535 8993
rect 45738 8956 45744 8968
rect 44192 8928 44312 8956
rect 45112 8928 45744 8956
rect 41322 8888 41328 8900
rect 41248 8860 41328 8888
rect 37976 8848 37982 8860
rect 41322 8848 41328 8860
rect 41380 8848 41386 8900
rect 44284 8888 44312 8928
rect 45738 8916 45744 8928
rect 45796 8956 45802 8968
rect 46201 8959 46259 8965
rect 46201 8956 46213 8959
rect 45796 8928 46213 8956
rect 45796 8916 45802 8928
rect 46201 8925 46213 8928
rect 46247 8925 46259 8959
rect 46934 8956 46940 8968
rect 46895 8928 46940 8956
rect 46201 8919 46259 8925
rect 46934 8916 46940 8928
rect 46992 8916 46998 8968
rect 47872 8956 47900 8996
rect 47946 8984 47952 9036
rect 48004 9024 48010 9036
rect 48004 8996 48049 9024
rect 48004 8984 48010 8996
rect 48682 8956 48688 8968
rect 47872 8928 48688 8956
rect 48682 8916 48688 8928
rect 48740 8916 48746 8968
rect 48792 8956 48820 9064
rect 49421 9061 49433 9095
rect 49467 9092 49479 9095
rect 50801 9095 50859 9101
rect 50801 9092 50813 9095
rect 49467 9064 50813 9092
rect 49467 9061 49479 9064
rect 49421 9055 49479 9061
rect 50801 9061 50813 9064
rect 50847 9061 50859 9095
rect 50801 9055 50859 9061
rect 49602 9024 49608 9036
rect 49563 8996 49608 9024
rect 49602 8984 49608 8996
rect 49660 8984 49666 9036
rect 49973 9027 50031 9033
rect 49973 8993 49985 9027
rect 50019 9024 50031 9027
rect 50430 9024 50436 9036
rect 50019 8996 50436 9024
rect 50019 8993 50031 8996
rect 49973 8987 50031 8993
rect 50430 8984 50436 8996
rect 50488 8984 50494 9036
rect 51442 9024 51448 9036
rect 51403 8996 51448 9024
rect 51442 8984 51448 8996
rect 51500 8984 51506 9036
rect 51718 8984 51724 9036
rect 51776 9024 51782 9036
rect 51920 9033 51948 9132
rect 56060 9132 58348 9160
rect 52914 9092 52920 9104
rect 52840 9064 52920 9092
rect 52840 9033 52868 9064
rect 52914 9052 52920 9064
rect 52972 9052 52978 9104
rect 54662 9092 54668 9104
rect 53024 9064 54668 9092
rect 51813 9027 51871 9033
rect 51813 9024 51825 9027
rect 51776 8996 51825 9024
rect 51776 8984 51782 8996
rect 51813 8993 51825 8996
rect 51859 8993 51871 9027
rect 51813 8987 51871 8993
rect 51905 9027 51963 9033
rect 51905 8993 51917 9027
rect 51951 8993 51963 9027
rect 52825 9027 52883 9033
rect 52825 9024 52837 9027
rect 51905 8987 51963 8993
rect 52104 8996 52837 9024
rect 51350 8956 51356 8968
rect 48792 8928 51212 8956
rect 51311 8928 51356 8956
rect 44284 8860 44588 8888
rect 34848 8792 37136 8820
rect 34848 8780 34854 8792
rect 37734 8780 37740 8832
rect 37792 8820 37798 8832
rect 40034 8820 40040 8832
rect 37792 8792 40040 8820
rect 37792 8780 37798 8792
rect 40034 8780 40040 8792
rect 40092 8780 40098 8832
rect 40129 8823 40187 8829
rect 40129 8789 40141 8823
rect 40175 8820 40187 8823
rect 44450 8820 44456 8832
rect 40175 8792 44456 8820
rect 40175 8789 40187 8792
rect 40129 8783 40187 8789
rect 44450 8780 44456 8792
rect 44508 8780 44514 8832
rect 44560 8820 44588 8860
rect 44818 8848 44824 8900
rect 44876 8888 44882 8900
rect 45097 8891 45155 8897
rect 45097 8888 45109 8891
rect 44876 8860 45109 8888
rect 44876 8848 44882 8860
rect 45097 8857 45109 8860
rect 45143 8857 45155 8891
rect 45097 8851 45155 8857
rect 47854 8848 47860 8900
rect 47912 8888 47918 8900
rect 49602 8888 49608 8900
rect 47912 8860 49608 8888
rect 47912 8848 47918 8860
rect 49602 8848 49608 8860
rect 49660 8848 49666 8900
rect 51184 8888 51212 8928
rect 51350 8916 51356 8928
rect 51408 8916 51414 8968
rect 52104 8888 52132 8996
rect 52825 8993 52837 8996
rect 52871 8993 52883 9027
rect 52825 8987 52883 8993
rect 53024 8965 53052 9064
rect 54662 9052 54668 9064
rect 54720 9052 54726 9104
rect 56060 9101 56088 9132
rect 58342 9120 58348 9132
rect 58400 9120 58406 9172
rect 56045 9095 56103 9101
rect 56045 9061 56057 9095
rect 56091 9061 56103 9095
rect 58066 9092 58072 9104
rect 58027 9064 58072 9092
rect 56045 9055 56103 9061
rect 58066 9052 58072 9064
rect 58124 9052 58130 9104
rect 58544 9064 59124 9092
rect 53650 8984 53656 9036
rect 53708 9024 53714 9036
rect 54754 9024 54760 9036
rect 53708 8996 54760 9024
rect 53708 8984 53714 8996
rect 54754 8984 54760 8996
rect 54812 8984 54818 9036
rect 54938 8984 54944 9036
rect 54996 9024 55002 9036
rect 56686 9024 56692 9036
rect 54996 8996 56692 9024
rect 54996 8984 55002 8996
rect 56686 8984 56692 8996
rect 56744 8984 56750 9036
rect 57054 9024 57060 9036
rect 57015 8996 57060 9024
rect 57054 8984 57060 8996
rect 57112 8984 57118 9036
rect 57238 9024 57244 9036
rect 57199 8996 57244 9024
rect 57238 8984 57244 8996
rect 57296 8984 57302 9036
rect 58544 9024 58572 9064
rect 58710 9024 58716 9036
rect 57992 8996 58572 9024
rect 58671 8996 58716 9024
rect 52972 8959 53052 8965
rect 52972 8925 52984 8959
rect 53018 8928 53052 8959
rect 53190 8956 53196 8968
rect 53151 8928 53196 8956
rect 53018 8925 53030 8928
rect 52972 8919 53030 8925
rect 53190 8916 53196 8928
rect 53248 8916 53254 8968
rect 54665 8959 54723 8965
rect 54665 8925 54677 8959
rect 54711 8956 54723 8959
rect 54846 8956 54852 8968
rect 54711 8928 54852 8956
rect 54711 8925 54723 8928
rect 54665 8919 54723 8925
rect 54846 8916 54852 8928
rect 54904 8916 54910 8968
rect 56781 8959 56839 8965
rect 56781 8925 56793 8959
rect 56827 8925 56839 8959
rect 57072 8956 57100 8984
rect 57992 8956 58020 8996
rect 58710 8984 58716 8996
rect 58768 8984 58774 9036
rect 59096 9033 59124 9064
rect 59081 9027 59139 9033
rect 59081 8993 59093 9027
rect 59127 9024 59139 9027
rect 59262 9024 59268 9036
rect 59127 8996 59268 9024
rect 59127 8993 59139 8996
rect 59081 8987 59139 8993
rect 59262 8984 59268 8996
rect 59320 8984 59326 9036
rect 60182 9024 60188 9036
rect 60143 8996 60188 9024
rect 60182 8984 60188 8996
rect 60240 8984 60246 9036
rect 60277 9027 60335 9033
rect 60277 8993 60289 9027
rect 60323 8993 60335 9027
rect 60277 8987 60335 8993
rect 58802 8956 58808 8968
rect 57072 8928 58020 8956
rect 58763 8928 58808 8956
rect 56781 8919 56839 8925
rect 51184 8860 52132 8888
rect 52178 8848 52184 8900
rect 52236 8888 52242 8900
rect 53285 8891 53343 8897
rect 53285 8888 53297 8891
rect 52236 8860 53297 8888
rect 52236 8848 52242 8860
rect 53285 8857 53297 8860
rect 53331 8857 53343 8891
rect 55030 8888 55036 8900
rect 53285 8851 53343 8857
rect 54864 8860 55036 8888
rect 45186 8820 45192 8832
rect 44560 8792 45192 8820
rect 45186 8780 45192 8792
rect 45244 8780 45250 8832
rect 45830 8780 45836 8832
rect 45888 8820 45894 8832
rect 47765 8823 47823 8829
rect 47765 8820 47777 8823
rect 45888 8792 47777 8820
rect 45888 8780 45894 8792
rect 47765 8789 47777 8792
rect 47811 8820 47823 8823
rect 49234 8820 49240 8832
rect 47811 8792 49240 8820
rect 47811 8789 47823 8792
rect 47765 8783 47823 8789
rect 49234 8780 49240 8792
rect 49292 8780 49298 8832
rect 49418 8780 49424 8832
rect 49476 8820 49482 8832
rect 53101 8823 53159 8829
rect 53101 8820 53113 8823
rect 49476 8792 53113 8820
rect 49476 8780 49482 8792
rect 53101 8789 53113 8792
rect 53147 8820 53159 8823
rect 54864 8820 54892 8860
rect 55030 8848 55036 8860
rect 55088 8848 55094 8900
rect 53147 8792 54892 8820
rect 54941 8823 54999 8829
rect 53147 8789 53159 8792
rect 53101 8783 53159 8789
rect 54941 8789 54953 8823
rect 54987 8820 54999 8823
rect 55306 8820 55312 8832
rect 54987 8792 55312 8820
rect 54987 8789 54999 8792
rect 54941 8783 54999 8789
rect 55306 8780 55312 8792
rect 55364 8780 55370 8832
rect 56796 8820 56824 8919
rect 58802 8916 58808 8928
rect 58860 8916 58866 8968
rect 59170 8956 59176 8968
rect 59131 8928 59176 8956
rect 59170 8916 59176 8928
rect 59228 8916 59234 8968
rect 56870 8848 56876 8900
rect 56928 8888 56934 8900
rect 60292 8888 60320 8987
rect 56928 8860 60320 8888
rect 56928 8848 56934 8860
rect 60461 8823 60519 8829
rect 60461 8820 60473 8823
rect 56796 8792 60473 8820
rect 60461 8789 60473 8792
rect 60507 8789 60519 8823
rect 60461 8783 60519 8789
rect 1104 8730 62192 8752
rect 1104 8678 11163 8730
rect 11215 8678 11227 8730
rect 11279 8678 11291 8730
rect 11343 8678 11355 8730
rect 11407 8678 31526 8730
rect 31578 8678 31590 8730
rect 31642 8678 31654 8730
rect 31706 8678 31718 8730
rect 31770 8678 51888 8730
rect 51940 8678 51952 8730
rect 52004 8678 52016 8730
rect 52068 8678 52080 8730
rect 52132 8678 62192 8730
rect 1104 8656 62192 8678
rect 1949 8619 2007 8625
rect 1949 8585 1961 8619
rect 1995 8616 2007 8619
rect 2774 8616 2780 8628
rect 1995 8588 2780 8616
rect 1995 8585 2007 8588
rect 1949 8579 2007 8585
rect 2774 8576 2780 8588
rect 2832 8576 2838 8628
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 4120 8588 4261 8616
rect 4120 8576 4126 8588
rect 4249 8585 4261 8588
rect 4295 8585 4307 8619
rect 4249 8579 4307 8585
rect 5537 8619 5595 8625
rect 5537 8585 5549 8619
rect 5583 8616 5595 8619
rect 5626 8616 5632 8628
rect 5583 8588 5632 8616
rect 5583 8585 5595 8588
rect 5537 8579 5595 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 9677 8619 9735 8625
rect 9677 8585 9689 8619
rect 9723 8616 9735 8619
rect 11514 8616 11520 8628
rect 9723 8588 11520 8616
rect 9723 8585 9735 8588
rect 9677 8579 9735 8585
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 14274 8616 14280 8628
rect 13372 8588 14280 8616
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8480 2927 8483
rect 3970 8480 3976 8492
rect 2915 8452 3976 8480
rect 2915 8449 2927 8452
rect 2869 8443 2927 8449
rect 3970 8440 3976 8452
rect 4028 8480 4034 8492
rect 8386 8480 8392 8492
rect 4028 8452 8156 8480
rect 8347 8452 8392 8480
rect 4028 8440 4034 8452
rect 1854 8412 1860 8424
rect 1815 8384 1860 8412
rect 1854 8372 1860 8384
rect 1912 8372 1918 8424
rect 3142 8412 3148 8424
rect 3103 8384 3148 8412
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 5350 8412 5356 8424
rect 5311 8384 5356 8412
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 8128 8421 8156 8452
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8480 12955 8483
rect 13372 8480 13400 8588
rect 14274 8576 14280 8588
rect 14332 8576 14338 8628
rect 19426 8576 19432 8628
rect 19484 8616 19490 8628
rect 21085 8619 21143 8625
rect 19484 8588 20852 8616
rect 19484 8576 19490 8588
rect 13538 8548 13544 8560
rect 13499 8520 13544 8548
rect 13538 8508 13544 8520
rect 13596 8508 13602 8560
rect 20714 8548 20720 8560
rect 14844 8520 20720 8548
rect 14737 8483 14795 8489
rect 14737 8480 14749 8483
rect 12943 8452 13400 8480
rect 13648 8452 14749 8480
rect 12943 8449 12955 8452
rect 12897 8443 12955 8449
rect 8113 8415 8171 8421
rect 8113 8381 8125 8415
rect 8159 8412 8171 8415
rect 8662 8412 8668 8424
rect 8159 8384 8668 8412
rect 8159 8381 8171 8384
rect 8113 8375 8171 8381
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 10042 8372 10048 8424
rect 10100 8412 10106 8424
rect 10597 8415 10655 8421
rect 10597 8412 10609 8415
rect 10100 8384 10609 8412
rect 10100 8372 10106 8384
rect 10597 8381 10609 8384
rect 10643 8381 10655 8415
rect 10597 8375 10655 8381
rect 10612 8276 10640 8375
rect 10870 8372 10876 8424
rect 10928 8412 10934 8424
rect 10965 8415 11023 8421
rect 10965 8412 10977 8415
rect 10928 8384 10977 8412
rect 10928 8372 10934 8384
rect 10965 8381 10977 8384
rect 11011 8381 11023 8415
rect 11146 8412 11152 8424
rect 11107 8384 11152 8412
rect 10965 8375 11023 8381
rect 11146 8372 11152 8384
rect 11204 8412 11210 8424
rect 11606 8412 11612 8424
rect 11204 8384 11612 8412
rect 11204 8372 11210 8384
rect 11606 8372 11612 8384
rect 11664 8372 11670 8424
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8381 13323 8415
rect 13265 8375 13323 8381
rect 13280 8344 13308 8375
rect 13354 8372 13360 8424
rect 13412 8412 13418 8424
rect 13648 8421 13676 8452
rect 14737 8449 14749 8452
rect 14783 8449 14795 8483
rect 14737 8443 14795 8449
rect 13633 8415 13691 8421
rect 13633 8412 13645 8415
rect 13412 8384 13645 8412
rect 13412 8372 13418 8384
rect 13633 8381 13645 8384
rect 13679 8381 13691 8415
rect 14642 8412 14648 8424
rect 14555 8384 14648 8412
rect 13633 8375 13691 8381
rect 14642 8372 14648 8384
rect 14700 8412 14706 8424
rect 14844 8412 14872 8520
rect 20714 8508 20720 8520
rect 20772 8508 20778 8560
rect 20824 8548 20852 8588
rect 21085 8585 21097 8619
rect 21131 8616 21143 8619
rect 21818 8616 21824 8628
rect 21131 8588 21824 8616
rect 21131 8585 21143 8588
rect 21085 8579 21143 8585
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 22002 8576 22008 8628
rect 22060 8616 22066 8628
rect 32030 8616 32036 8628
rect 22060 8588 32036 8616
rect 22060 8576 22066 8588
rect 32030 8576 32036 8588
rect 32088 8616 32094 8628
rect 33042 8616 33048 8628
rect 32088 8588 33048 8616
rect 32088 8576 32094 8588
rect 33042 8576 33048 8588
rect 33100 8576 33106 8628
rect 34054 8576 34060 8628
rect 34112 8616 34118 8628
rect 34112 8588 34652 8616
rect 34112 8576 34118 8588
rect 22186 8548 22192 8560
rect 20824 8520 22192 8548
rect 22186 8508 22192 8520
rect 22244 8508 22250 8560
rect 22370 8508 22376 8560
rect 22428 8548 22434 8560
rect 22428 8520 22692 8548
rect 22428 8508 22434 8520
rect 15562 8440 15568 8492
rect 15620 8480 15626 8492
rect 15933 8483 15991 8489
rect 15933 8480 15945 8483
rect 15620 8452 15945 8480
rect 15620 8440 15626 8452
rect 15933 8449 15945 8452
rect 15979 8480 15991 8483
rect 20162 8480 20168 8492
rect 15979 8452 20168 8480
rect 15979 8449 15991 8452
rect 15933 8443 15991 8449
rect 20162 8440 20168 8452
rect 20220 8440 20226 8492
rect 21008 8452 22416 8480
rect 16022 8412 16028 8424
rect 14700 8384 14872 8412
rect 15983 8384 16028 8412
rect 14700 8372 14706 8384
rect 16022 8372 16028 8384
rect 16080 8412 16086 8424
rect 18506 8412 18512 8424
rect 16080 8384 18512 8412
rect 16080 8372 16086 8384
rect 18506 8372 18512 8384
rect 18564 8372 18570 8424
rect 18690 8412 18696 8424
rect 18651 8384 18696 8412
rect 18690 8372 18696 8384
rect 18748 8372 18754 8424
rect 19061 8415 19119 8421
rect 19061 8381 19073 8415
rect 19107 8412 19119 8415
rect 19889 8415 19947 8421
rect 19889 8412 19901 8415
rect 19107 8384 19901 8412
rect 19107 8381 19119 8384
rect 19061 8375 19119 8381
rect 19889 8381 19901 8384
rect 19935 8381 19947 8415
rect 20070 8412 20076 8424
rect 20031 8384 20076 8412
rect 19889 8375 19947 8381
rect 16485 8347 16543 8353
rect 16485 8344 16497 8347
rect 13280 8316 16497 8344
rect 16485 8313 16497 8316
rect 16531 8344 16543 8347
rect 17586 8344 17592 8356
rect 16531 8316 17592 8344
rect 16531 8313 16543 8316
rect 16485 8307 16543 8313
rect 17586 8304 17592 8316
rect 17644 8304 17650 8356
rect 19904 8344 19932 8375
rect 20070 8372 20076 8384
rect 20128 8372 20134 8424
rect 20530 8412 20536 8424
rect 20491 8384 20536 8412
rect 20530 8372 20536 8384
rect 20588 8372 20594 8424
rect 20622 8372 20628 8424
rect 20680 8412 20686 8424
rect 20680 8384 20725 8412
rect 20680 8372 20686 8384
rect 20806 8372 20812 8424
rect 20864 8412 20870 8424
rect 21008 8412 21036 8452
rect 20864 8384 21036 8412
rect 20864 8372 20870 8384
rect 22186 8372 22192 8424
rect 22244 8412 22250 8424
rect 22281 8415 22339 8421
rect 22281 8412 22293 8415
rect 22244 8384 22293 8412
rect 22244 8372 22250 8384
rect 22281 8381 22293 8384
rect 22327 8381 22339 8415
rect 22281 8375 22339 8381
rect 20898 8344 20904 8356
rect 19904 8316 20904 8344
rect 20898 8304 20904 8316
rect 20956 8304 20962 8356
rect 21818 8304 21824 8356
rect 21876 8344 21882 8356
rect 22097 8347 22155 8353
rect 22097 8344 22109 8347
rect 21876 8316 22109 8344
rect 21876 8304 21882 8316
rect 22097 8313 22109 8316
rect 22143 8313 22155 8347
rect 22388 8344 22416 8452
rect 22462 8440 22468 8492
rect 22520 8480 22526 8492
rect 22557 8483 22615 8489
rect 22557 8480 22569 8483
rect 22520 8452 22569 8480
rect 22520 8440 22526 8452
rect 22557 8449 22569 8452
rect 22603 8449 22615 8483
rect 22664 8480 22692 8520
rect 23842 8508 23848 8560
rect 23900 8548 23906 8560
rect 30834 8548 30840 8560
rect 23900 8520 23945 8548
rect 24136 8520 30840 8548
rect 23900 8508 23906 8520
rect 24136 8480 24164 8520
rect 30834 8508 30840 8520
rect 30892 8548 30898 8560
rect 34624 8548 34652 8588
rect 36078 8576 36084 8628
rect 36136 8616 36142 8628
rect 37093 8619 37151 8625
rect 37093 8616 37105 8619
rect 36136 8588 37105 8616
rect 36136 8576 36142 8588
rect 37093 8585 37105 8588
rect 37139 8585 37151 8619
rect 37093 8579 37151 8585
rect 38381 8619 38439 8625
rect 38381 8585 38393 8619
rect 38427 8616 38439 8619
rect 39298 8616 39304 8628
rect 38427 8588 39304 8616
rect 38427 8585 38439 8588
rect 38381 8579 38439 8585
rect 39298 8576 39304 8588
rect 39356 8576 39362 8628
rect 39482 8616 39488 8628
rect 39443 8588 39488 8616
rect 39482 8576 39488 8588
rect 39540 8576 39546 8628
rect 41693 8619 41751 8625
rect 41693 8585 41705 8619
rect 41739 8616 41751 8619
rect 42058 8616 42064 8628
rect 41739 8588 42064 8616
rect 41739 8585 41751 8588
rect 41693 8579 41751 8585
rect 42058 8576 42064 8588
rect 42116 8576 42122 8628
rect 43717 8619 43775 8625
rect 43717 8585 43729 8619
rect 43763 8616 43775 8619
rect 44634 8616 44640 8628
rect 43763 8588 44640 8616
rect 43763 8585 43775 8588
rect 43717 8579 43775 8585
rect 44634 8576 44640 8588
rect 44692 8576 44698 8628
rect 48130 8576 48136 8628
rect 48188 8616 48194 8628
rect 50338 8616 50344 8628
rect 48188 8588 50344 8616
rect 48188 8576 48194 8588
rect 50338 8576 50344 8588
rect 50396 8576 50402 8628
rect 50430 8576 50436 8628
rect 50488 8616 50494 8628
rect 50525 8619 50583 8625
rect 50525 8616 50537 8619
rect 50488 8588 50537 8616
rect 50488 8576 50494 8588
rect 50525 8585 50537 8588
rect 50571 8585 50583 8619
rect 52730 8616 52736 8628
rect 52691 8588 52736 8616
rect 50525 8579 50583 8585
rect 52730 8576 52736 8588
rect 52788 8576 52794 8628
rect 55030 8576 55036 8628
rect 55088 8616 55094 8628
rect 58526 8616 58532 8628
rect 55088 8588 58532 8616
rect 55088 8576 55094 8588
rect 58526 8576 58532 8588
rect 58584 8576 58590 8628
rect 36538 8548 36544 8560
rect 30892 8520 34560 8548
rect 34624 8520 36544 8548
rect 30892 8508 30898 8520
rect 34532 8492 34560 8520
rect 36538 8508 36544 8520
rect 36596 8508 36602 8560
rect 36998 8508 37004 8560
rect 37056 8548 37062 8560
rect 42150 8548 42156 8560
rect 37056 8520 42156 8548
rect 37056 8508 37062 8520
rect 42150 8508 42156 8520
rect 42208 8508 42214 8560
rect 42334 8508 42340 8560
rect 42392 8548 42398 8560
rect 42794 8548 42800 8560
rect 42392 8520 42800 8548
rect 42392 8508 42398 8520
rect 25685 8483 25743 8489
rect 22664 8452 24164 8480
rect 25240 8452 25544 8480
rect 22557 8443 22615 8449
rect 23382 8372 23388 8424
rect 23440 8412 23446 8424
rect 23661 8415 23719 8421
rect 23661 8412 23673 8415
rect 23440 8384 23673 8412
rect 23440 8372 23446 8384
rect 23661 8381 23673 8384
rect 23707 8381 23719 8415
rect 23661 8375 23719 8381
rect 24854 8372 24860 8424
rect 24912 8412 24918 8424
rect 25240 8421 25268 8452
rect 25225 8415 25283 8421
rect 25225 8412 25237 8415
rect 24912 8384 25237 8412
rect 24912 8372 24918 8384
rect 25225 8381 25237 8384
rect 25271 8381 25283 8415
rect 25406 8412 25412 8424
rect 25367 8384 25412 8412
rect 25225 8375 25283 8381
rect 25406 8372 25412 8384
rect 25464 8372 25470 8424
rect 25516 8412 25544 8452
rect 25685 8449 25697 8483
rect 25731 8480 25743 8483
rect 26510 8480 26516 8492
rect 25731 8452 26516 8480
rect 25731 8449 25743 8452
rect 25685 8443 25743 8449
rect 26510 8440 26516 8452
rect 26568 8440 26574 8492
rect 26697 8483 26755 8489
rect 26697 8449 26709 8483
rect 26743 8480 26755 8483
rect 27798 8480 27804 8492
rect 26743 8452 27804 8480
rect 26743 8449 26755 8452
rect 26697 8443 26755 8449
rect 27798 8440 27804 8452
rect 27856 8440 27862 8492
rect 30193 8483 30251 8489
rect 30193 8449 30205 8483
rect 30239 8480 30251 8483
rect 30374 8480 30380 8492
rect 30239 8452 30380 8480
rect 30239 8449 30251 8452
rect 30193 8443 30251 8449
rect 30374 8440 30380 8452
rect 30432 8440 30438 8492
rect 31846 8480 31852 8492
rect 31807 8452 31852 8480
rect 31846 8440 31852 8452
rect 31904 8440 31910 8492
rect 32401 8483 32459 8489
rect 32401 8449 32413 8483
rect 32447 8480 32459 8483
rect 33134 8480 33140 8492
rect 32447 8452 33140 8480
rect 32447 8449 32459 8452
rect 32401 8443 32459 8449
rect 33134 8440 33140 8452
rect 33192 8440 33198 8492
rect 33597 8483 33655 8489
rect 33597 8449 33609 8483
rect 33643 8480 33655 8483
rect 33870 8480 33876 8492
rect 33643 8452 33876 8480
rect 33643 8449 33655 8452
rect 33597 8443 33655 8449
rect 33870 8440 33876 8452
rect 33928 8440 33934 8492
rect 34514 8440 34520 8492
rect 34572 8480 34578 8492
rect 34572 8452 42288 8480
rect 34572 8440 34578 8452
rect 26878 8412 26884 8424
rect 25516 8384 26884 8412
rect 26878 8372 26884 8384
rect 26936 8372 26942 8424
rect 26973 8415 27031 8421
rect 26973 8381 26985 8415
rect 27019 8381 27031 8415
rect 26973 8375 27031 8381
rect 26988 8344 27016 8375
rect 27062 8372 27068 8424
rect 27120 8412 27126 8424
rect 27341 8415 27399 8421
rect 27341 8412 27353 8415
rect 27120 8384 27353 8412
rect 27120 8372 27126 8384
rect 27341 8381 27353 8384
rect 27387 8412 27399 8415
rect 27387 8384 27752 8412
rect 27387 8381 27399 8384
rect 27341 8375 27399 8381
rect 27430 8344 27436 8356
rect 22388 8316 27436 8344
rect 22097 8307 22155 8313
rect 27430 8304 27436 8316
rect 27488 8304 27494 8356
rect 27614 8344 27620 8356
rect 27575 8316 27620 8344
rect 27614 8304 27620 8316
rect 27672 8304 27678 8356
rect 27724 8344 27752 8384
rect 29546 8372 29552 8424
rect 29604 8412 29610 8424
rect 29641 8415 29699 8421
rect 29641 8412 29653 8415
rect 29604 8384 29653 8412
rect 29604 8372 29610 8384
rect 29641 8381 29653 8384
rect 29687 8381 29699 8415
rect 29641 8375 29699 8381
rect 29730 8372 29736 8424
rect 29788 8412 29794 8424
rect 31018 8412 31024 8424
rect 29788 8384 31024 8412
rect 29788 8372 29794 8384
rect 31018 8372 31024 8384
rect 31076 8372 31082 8424
rect 31941 8415 31999 8421
rect 31941 8381 31953 8415
rect 31987 8412 31999 8415
rect 32306 8412 32312 8424
rect 31987 8384 32312 8412
rect 31987 8381 31999 8384
rect 31941 8375 31999 8381
rect 32306 8372 32312 8384
rect 32364 8372 32370 8424
rect 33226 8412 33232 8424
rect 33187 8384 33232 8412
rect 33226 8372 33232 8384
rect 33284 8372 33290 8424
rect 33778 8412 33784 8424
rect 33739 8384 33784 8412
rect 33778 8372 33784 8384
rect 33836 8372 33842 8424
rect 34882 8412 34888 8424
rect 34843 8384 34888 8412
rect 34882 8372 34888 8384
rect 34940 8372 34946 8424
rect 35434 8412 35440 8424
rect 35395 8384 35440 8412
rect 35434 8372 35440 8384
rect 35492 8372 35498 8424
rect 35710 8412 35716 8424
rect 35544 8384 35716 8412
rect 35544 8344 35572 8384
rect 35710 8372 35716 8384
rect 35768 8372 35774 8424
rect 36814 8412 36820 8424
rect 35820 8384 36308 8412
rect 36775 8384 36820 8412
rect 27724 8316 35572 8344
rect 35618 8304 35624 8356
rect 35676 8344 35682 8356
rect 35820 8344 35848 8384
rect 35676 8316 35848 8344
rect 35989 8347 36047 8353
rect 35676 8304 35682 8316
rect 35989 8313 36001 8347
rect 36035 8344 36047 8347
rect 36170 8344 36176 8356
rect 36035 8316 36176 8344
rect 36035 8313 36047 8316
rect 35989 8307 36047 8313
rect 36170 8304 36176 8316
rect 36228 8304 36234 8356
rect 36280 8344 36308 8384
rect 36814 8372 36820 8384
rect 36872 8372 36878 8424
rect 36909 8415 36967 8421
rect 36909 8381 36921 8415
rect 36955 8412 36967 8415
rect 37274 8412 37280 8424
rect 36955 8384 37280 8412
rect 36955 8381 36967 8384
rect 36909 8375 36967 8381
rect 37274 8372 37280 8384
rect 37332 8412 37338 8424
rect 38197 8415 38255 8421
rect 38197 8412 38209 8415
rect 37332 8384 38209 8412
rect 37332 8372 37338 8384
rect 38197 8381 38209 8384
rect 38243 8381 38255 8415
rect 38197 8375 38255 8381
rect 38286 8372 38292 8424
rect 38344 8412 38350 8424
rect 39301 8415 39359 8421
rect 39301 8412 39313 8415
rect 38344 8384 39313 8412
rect 38344 8372 38350 8384
rect 39301 8381 39313 8384
rect 39347 8381 39359 8415
rect 39301 8375 39359 8381
rect 40034 8372 40040 8424
rect 40092 8412 40098 8424
rect 40497 8415 40555 8421
rect 40497 8412 40509 8415
rect 40092 8384 40509 8412
rect 40092 8372 40098 8384
rect 40497 8381 40509 8384
rect 40543 8412 40555 8415
rect 41414 8412 41420 8424
rect 40543 8384 41420 8412
rect 40543 8381 40555 8384
rect 40497 8375 40555 8381
rect 41414 8372 41420 8384
rect 41472 8372 41478 8424
rect 42150 8372 42156 8424
rect 42208 8412 42214 8424
rect 42260 8421 42288 8452
rect 42245 8415 42303 8421
rect 42245 8412 42257 8415
rect 42208 8384 42257 8412
rect 42208 8372 42214 8384
rect 42245 8381 42257 8384
rect 42291 8381 42303 8415
rect 42245 8375 42303 8381
rect 42337 8415 42395 8421
rect 42337 8381 42349 8415
rect 42383 8412 42395 8415
rect 42426 8412 42432 8424
rect 42383 8384 42432 8412
rect 42383 8381 42395 8384
rect 42337 8375 42395 8381
rect 42426 8372 42432 8384
rect 42484 8372 42490 8424
rect 42628 8421 42656 8520
rect 42794 8508 42800 8520
rect 42852 8508 42858 8560
rect 46201 8551 46259 8557
rect 46201 8517 46213 8551
rect 46247 8517 46259 8551
rect 46201 8511 46259 8517
rect 46216 8480 46244 8511
rect 46290 8508 46296 8560
rect 46348 8548 46354 8560
rect 46348 8520 48228 8548
rect 46348 8508 46354 8520
rect 46934 8480 46940 8492
rect 42720 8452 46244 8480
rect 46895 8452 46940 8480
rect 42613 8415 42671 8421
rect 42613 8381 42625 8415
rect 42659 8381 42671 8415
rect 42613 8375 42671 8381
rect 42720 8344 42748 8452
rect 46934 8440 46940 8452
rect 46992 8440 46998 8492
rect 42797 8415 42855 8421
rect 42797 8381 42809 8415
rect 42843 8412 42855 8415
rect 42886 8412 42892 8424
rect 42843 8384 42892 8412
rect 42843 8381 42855 8384
rect 42797 8375 42855 8381
rect 42886 8372 42892 8384
rect 42944 8372 42950 8424
rect 44174 8372 44180 8424
rect 44232 8421 44238 8424
rect 44232 8415 44249 8421
rect 44237 8381 44249 8415
rect 44358 8412 44364 8424
rect 44319 8384 44364 8412
rect 44232 8375 44249 8381
rect 44232 8372 44238 8375
rect 44358 8372 44364 8384
rect 44416 8372 44422 8424
rect 44450 8372 44456 8424
rect 44508 8412 44514 8424
rect 44637 8415 44695 8421
rect 44637 8412 44649 8415
rect 44508 8384 44649 8412
rect 44508 8372 44514 8384
rect 44637 8381 44649 8384
rect 44683 8381 44695 8415
rect 44818 8412 44824 8424
rect 44779 8384 44824 8412
rect 44637 8375 44695 8381
rect 44818 8372 44824 8384
rect 44876 8372 44882 8424
rect 45830 8412 45836 8424
rect 45791 8384 45836 8412
rect 45830 8372 45836 8384
rect 45888 8372 45894 8424
rect 46290 8412 46296 8424
rect 46251 8384 46296 8412
rect 46290 8372 46296 8384
rect 46348 8372 46354 8424
rect 46842 8412 46848 8424
rect 46803 8384 46848 8412
rect 46842 8372 46848 8384
rect 46900 8372 46906 8424
rect 48200 8421 48228 8520
rect 51350 8508 51356 8560
rect 51408 8548 51414 8560
rect 55214 8548 55220 8560
rect 51408 8520 55220 8548
rect 51408 8508 51414 8520
rect 48406 8440 48412 8492
rect 48464 8480 48470 8492
rect 53285 8483 53343 8489
rect 53285 8480 53297 8483
rect 48464 8452 53297 8480
rect 48464 8440 48470 8452
rect 53285 8449 53297 8452
rect 53331 8449 53343 8483
rect 54938 8480 54944 8492
rect 53285 8443 53343 8449
rect 53576 8452 54944 8480
rect 48200 8415 48283 8421
rect 48200 8384 48237 8415
rect 48225 8381 48237 8384
rect 48271 8381 48283 8415
rect 50246 8412 50252 8424
rect 50207 8384 50252 8412
rect 48225 8375 48283 8381
rect 50246 8372 50252 8384
rect 50304 8372 50310 8424
rect 50338 8372 50344 8424
rect 50396 8412 50402 8424
rect 52178 8412 52184 8424
rect 50396 8384 52184 8412
rect 50396 8372 50402 8384
rect 52178 8372 52184 8384
rect 52236 8372 52242 8424
rect 53190 8412 53196 8424
rect 53248 8421 53254 8424
rect 53248 8415 53265 8421
rect 53117 8384 53196 8412
rect 53190 8372 53196 8384
rect 53253 8412 53265 8415
rect 53576 8412 53604 8452
rect 54938 8440 54944 8452
rect 54996 8440 55002 8492
rect 55048 8489 55076 8520
rect 55214 8508 55220 8520
rect 55272 8508 55278 8560
rect 58802 8548 58808 8560
rect 58763 8520 58808 8548
rect 58802 8508 58808 8520
rect 58860 8508 58866 8560
rect 55033 8483 55091 8489
rect 55033 8449 55045 8483
rect 55079 8449 55091 8483
rect 55033 8443 55091 8449
rect 55125 8483 55183 8489
rect 55125 8449 55137 8483
rect 55171 8480 55183 8483
rect 59170 8480 59176 8492
rect 55171 8452 59176 8480
rect 55171 8449 55183 8452
rect 55125 8443 55183 8449
rect 59170 8440 59176 8452
rect 59228 8440 59234 8492
rect 53253 8384 53604 8412
rect 53253 8381 53265 8384
rect 53248 8375 53265 8381
rect 53248 8372 53254 8375
rect 53650 8372 53656 8424
rect 53708 8412 53714 8424
rect 53837 8415 53895 8421
rect 53708 8384 53753 8412
rect 53708 8372 53714 8384
rect 53837 8381 53849 8415
rect 53883 8381 53895 8415
rect 55858 8412 55864 8424
rect 55819 8384 55864 8412
rect 53837 8375 53895 8381
rect 36280 8316 42748 8344
rect 46106 8304 46112 8356
rect 46164 8344 46170 8356
rect 47946 8344 47952 8356
rect 46164 8316 47952 8344
rect 46164 8304 46170 8316
rect 47946 8304 47952 8316
rect 48004 8344 48010 8356
rect 48041 8347 48099 8353
rect 48041 8344 48053 8347
rect 48004 8316 48053 8344
rect 48004 8304 48010 8316
rect 48041 8313 48053 8316
rect 48087 8313 48099 8347
rect 53852 8344 53880 8375
rect 55858 8372 55864 8384
rect 55916 8372 55922 8424
rect 55999 8415 56057 8421
rect 55999 8381 56011 8415
rect 56045 8412 56057 8415
rect 56318 8412 56324 8424
rect 56045 8384 56324 8412
rect 56045 8381 56057 8384
rect 55999 8375 56057 8381
rect 56318 8372 56324 8384
rect 56376 8372 56382 8424
rect 58526 8412 58532 8424
rect 58487 8384 58532 8412
rect 58526 8372 58532 8384
rect 58584 8372 58590 8424
rect 59262 8412 59268 8424
rect 59223 8384 59268 8412
rect 59262 8372 59268 8384
rect 59320 8372 59326 8424
rect 59541 8415 59599 8421
rect 59541 8381 59553 8415
rect 59587 8381 59599 8415
rect 59541 8375 59599 8381
rect 56870 8344 56876 8356
rect 48041 8307 48099 8313
rect 48148 8316 48360 8344
rect 19978 8276 19984 8288
rect 10612 8248 19984 8276
rect 19978 8236 19984 8248
rect 20036 8236 20042 8288
rect 20070 8236 20076 8288
rect 20128 8276 20134 8288
rect 30650 8276 30656 8288
rect 20128 8248 30656 8276
rect 20128 8236 20134 8248
rect 30650 8236 30656 8248
rect 30708 8236 30714 8288
rect 32766 8236 32772 8288
rect 32824 8276 32830 8288
rect 39758 8276 39764 8288
rect 32824 8248 39764 8276
rect 32824 8236 32830 8248
rect 39758 8236 39764 8248
rect 39816 8236 39822 8288
rect 40678 8276 40684 8288
rect 40591 8248 40684 8276
rect 40678 8236 40684 8248
rect 40736 8276 40742 8288
rect 44818 8276 44824 8288
rect 40736 8248 44824 8276
rect 40736 8236 40742 8248
rect 44818 8236 44824 8248
rect 44876 8236 44882 8288
rect 45554 8236 45560 8288
rect 45612 8276 45618 8288
rect 45649 8279 45707 8285
rect 45649 8276 45661 8279
rect 45612 8248 45661 8276
rect 45612 8236 45618 8248
rect 45649 8245 45661 8248
rect 45695 8276 45707 8279
rect 46014 8276 46020 8288
rect 45695 8248 46020 8276
rect 45695 8245 45707 8248
rect 45649 8239 45707 8245
rect 46014 8236 46020 8248
rect 46072 8236 46078 8288
rect 46382 8236 46388 8288
rect 46440 8276 46446 8288
rect 48148 8276 48176 8316
rect 48332 8285 48360 8316
rect 53852 8316 56876 8344
rect 46440 8248 48176 8276
rect 48317 8279 48375 8285
rect 46440 8236 46446 8248
rect 48317 8245 48329 8279
rect 48363 8245 48375 8279
rect 48317 8239 48375 8245
rect 49602 8236 49608 8288
rect 49660 8276 49666 8288
rect 50798 8276 50804 8288
rect 49660 8248 50804 8276
rect 49660 8236 49666 8248
rect 50798 8236 50804 8248
rect 50856 8276 50862 8288
rect 53852 8276 53880 8316
rect 56870 8304 56876 8316
rect 56928 8304 56934 8356
rect 56962 8304 56968 8356
rect 57020 8344 57026 8356
rect 59556 8344 59584 8375
rect 57020 8316 59584 8344
rect 57020 8304 57026 8316
rect 50856 8248 53880 8276
rect 50856 8236 50862 8248
rect 1104 8186 62192 8208
rect 1104 8134 21344 8186
rect 21396 8134 21408 8186
rect 21460 8134 21472 8186
rect 21524 8134 21536 8186
rect 21588 8134 41707 8186
rect 41759 8134 41771 8186
rect 41823 8134 41835 8186
rect 41887 8134 41899 8186
rect 41951 8134 62192 8186
rect 1104 8112 62192 8134
rect 9953 8075 10011 8081
rect 9953 8041 9965 8075
rect 9999 8072 10011 8075
rect 10778 8072 10784 8084
rect 9999 8044 10784 8072
rect 9999 8041 10011 8044
rect 9953 8035 10011 8041
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 15930 8072 15936 8084
rect 11992 8044 15936 8072
rect 4062 8004 4068 8016
rect 2976 7976 4068 8004
rect 2593 7939 2651 7945
rect 2593 7905 2605 7939
rect 2639 7936 2651 7939
rect 2866 7936 2872 7948
rect 2639 7908 2872 7936
rect 2639 7905 2651 7908
rect 2593 7899 2651 7905
rect 2866 7896 2872 7908
rect 2924 7896 2930 7948
rect 2976 7945 3004 7976
rect 4062 7964 4068 7976
rect 4120 7964 4126 8016
rect 4249 8007 4307 8013
rect 4249 7973 4261 8007
rect 4295 8004 4307 8007
rect 4338 8004 4344 8016
rect 4295 7976 4344 8004
rect 4295 7973 4307 7976
rect 4249 7967 4307 7973
rect 4338 7964 4344 7976
rect 4396 7964 4402 8016
rect 8205 8007 8263 8013
rect 8205 7973 8217 8007
rect 8251 8004 8263 8007
rect 11146 8004 11152 8016
rect 8251 7976 11152 8004
rect 8251 7973 8263 7976
rect 8205 7967 8263 7973
rect 11146 7964 11152 7976
rect 11204 7964 11210 8016
rect 2961 7939 3019 7945
rect 2961 7905 2973 7939
rect 3007 7905 3019 7939
rect 2961 7899 3019 7905
rect 3234 7896 3240 7948
rect 3292 7936 3298 7948
rect 4709 7939 4767 7945
rect 4709 7936 4721 7939
rect 3292 7908 4721 7936
rect 3292 7896 3298 7908
rect 4709 7905 4721 7908
rect 4755 7905 4767 7939
rect 5074 7936 5080 7948
rect 5035 7908 5080 7936
rect 4709 7899 4767 7905
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7936 5227 7939
rect 5626 7936 5632 7948
rect 5215 7908 5632 7936
rect 5215 7905 5227 7908
rect 5169 7899 5227 7905
rect 3050 7868 3056 7880
rect 2963 7840 3056 7868
rect 3050 7828 3056 7840
rect 3108 7868 3114 7880
rect 5184 7868 5212 7899
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 8389 7939 8447 7945
rect 8389 7936 8401 7939
rect 8352 7908 8401 7936
rect 8352 7896 8358 7908
rect 8389 7905 8401 7908
rect 8435 7905 8447 7939
rect 10318 7936 10324 7948
rect 10279 7908 10324 7936
rect 8389 7899 8447 7905
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 10686 7936 10692 7948
rect 10647 7908 10692 7936
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 11992 7945 12020 8044
rect 15930 8032 15936 8044
rect 15988 8032 15994 8084
rect 16482 8032 16488 8084
rect 16540 8072 16546 8084
rect 17678 8072 17684 8084
rect 16540 8044 17684 8072
rect 16540 8032 16546 8044
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 19702 8032 19708 8084
rect 19760 8072 19766 8084
rect 22094 8072 22100 8084
rect 19760 8044 22100 8072
rect 19760 8032 19766 8044
rect 22094 8032 22100 8044
rect 22152 8032 22158 8084
rect 22186 8032 22192 8084
rect 22244 8072 22250 8084
rect 22244 8044 30604 8072
rect 22244 8032 22250 8044
rect 12069 8007 12127 8013
rect 12069 7973 12081 8007
rect 12115 8004 12127 8007
rect 12710 8004 12716 8016
rect 12115 7976 12716 8004
rect 12115 7973 12127 7976
rect 12069 7967 12127 7973
rect 12710 7964 12716 7976
rect 12768 7964 12774 8016
rect 12820 7976 13952 8004
rect 10873 7939 10931 7945
rect 10873 7905 10885 7939
rect 10919 7905 10931 7939
rect 10873 7899 10931 7905
rect 11977 7939 12035 7945
rect 11977 7905 11989 7939
rect 12023 7905 12035 7939
rect 11977 7899 12035 7905
rect 12529 7939 12587 7945
rect 12529 7905 12541 7939
rect 12575 7936 12587 7939
rect 12618 7936 12624 7948
rect 12575 7908 12624 7936
rect 12575 7905 12587 7908
rect 12529 7899 12587 7905
rect 8754 7868 8760 7880
rect 3108 7840 5212 7868
rect 8715 7840 8760 7868
rect 3108 7828 3114 7840
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 10226 7868 10232 7880
rect 10187 7840 10232 7868
rect 10226 7828 10232 7840
rect 10284 7828 10290 7880
rect 10888 7868 10916 7899
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 12820 7868 12848 7976
rect 12897 7939 12955 7945
rect 12897 7905 12909 7939
rect 12943 7936 12955 7939
rect 13538 7936 13544 7948
rect 12943 7908 13544 7936
rect 12943 7905 12955 7908
rect 12897 7899 12955 7905
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 10888 7840 12848 7868
rect 12989 7871 13047 7877
rect 12989 7837 13001 7871
rect 13035 7868 13047 7871
rect 13814 7868 13820 7880
rect 13035 7840 13820 7868
rect 13035 7837 13047 7840
rect 12989 7831 13047 7837
rect 13814 7828 13820 7840
rect 13872 7828 13878 7880
rect 13924 7868 13952 7976
rect 14108 7976 17816 8004
rect 14108 7945 14136 7976
rect 14093 7939 14151 7945
rect 14093 7905 14105 7939
rect 14139 7905 14151 7939
rect 14093 7899 14151 7905
rect 14642 7896 14648 7948
rect 14700 7936 14706 7948
rect 15381 7939 15439 7945
rect 15381 7936 15393 7939
rect 14700 7908 15393 7936
rect 14700 7896 14706 7908
rect 15381 7905 15393 7908
rect 15427 7936 15439 7939
rect 16114 7936 16120 7948
rect 15427 7908 16120 7936
rect 15427 7905 15439 7908
rect 15381 7899 15439 7905
rect 16114 7896 16120 7908
rect 16172 7896 16178 7948
rect 17586 7936 17592 7948
rect 17547 7908 17592 7936
rect 17586 7896 17592 7908
rect 17644 7896 17650 7948
rect 17788 7945 17816 7976
rect 17862 7964 17868 8016
rect 17920 8004 17926 8016
rect 20438 8004 20444 8016
rect 17920 7976 20444 8004
rect 17920 7964 17926 7976
rect 20438 7964 20444 7976
rect 20496 7964 20502 8016
rect 20530 7964 20536 8016
rect 20588 8004 20594 8016
rect 26789 8007 26847 8013
rect 20588 7976 23796 8004
rect 20588 7964 20594 7976
rect 17773 7939 17831 7945
rect 17773 7905 17785 7939
rect 17819 7936 17831 7939
rect 19518 7936 19524 7948
rect 17819 7908 19435 7936
rect 19479 7908 19524 7936
rect 17819 7905 17831 7908
rect 17773 7899 17831 7905
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 13924 7840 15301 7868
rect 15289 7837 15301 7840
rect 15335 7868 15347 7871
rect 15838 7868 15844 7880
rect 15335 7840 15844 7868
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 16761 7871 16819 7877
rect 16761 7868 16773 7871
rect 16632 7840 16773 7868
rect 16632 7828 16638 7840
rect 16761 7837 16773 7840
rect 16807 7837 16819 7871
rect 16761 7831 16819 7837
rect 17313 7871 17371 7877
rect 17313 7837 17325 7871
rect 17359 7868 17371 7871
rect 18046 7868 18052 7880
rect 17359 7840 18052 7868
rect 17359 7837 17371 7840
rect 17313 7831 17371 7837
rect 18046 7828 18052 7840
rect 18104 7868 18110 7880
rect 18690 7868 18696 7880
rect 18104 7840 18696 7868
rect 18104 7828 18110 7840
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 18969 7871 19027 7877
rect 18969 7837 18981 7871
rect 19015 7868 19027 7871
rect 19242 7868 19248 7880
rect 19015 7840 19248 7868
rect 19015 7837 19027 7840
rect 18969 7831 19027 7837
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 19407 7868 19435 7908
rect 19518 7896 19524 7908
rect 19576 7896 19582 7948
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7936 19855 7939
rect 20622 7936 20628 7948
rect 19843 7908 20628 7936
rect 19843 7905 19855 7908
rect 19797 7899 19855 7905
rect 20622 7896 20628 7908
rect 20680 7896 20686 7948
rect 20806 7896 20812 7948
rect 20864 7936 20870 7948
rect 20901 7939 20959 7945
rect 20901 7936 20913 7939
rect 20864 7908 20913 7936
rect 20864 7896 20870 7908
rect 20901 7905 20913 7908
rect 20947 7905 20959 7939
rect 21082 7936 21088 7948
rect 20995 7908 21088 7936
rect 20901 7899 20959 7905
rect 21082 7896 21088 7908
rect 21140 7936 21146 7948
rect 22186 7936 22192 7948
rect 21140 7908 22192 7936
rect 21140 7896 21146 7908
rect 22186 7896 22192 7908
rect 22244 7896 22250 7948
rect 22465 7939 22523 7945
rect 22465 7905 22477 7939
rect 22511 7936 22523 7939
rect 22554 7936 22560 7948
rect 22511 7908 22560 7936
rect 22511 7905 22523 7908
rect 22465 7899 22523 7905
rect 22554 7896 22560 7908
rect 22612 7896 22618 7948
rect 23017 7939 23075 7945
rect 23017 7905 23029 7939
rect 23063 7936 23075 7939
rect 23658 7936 23664 7948
rect 23063 7908 23664 7936
rect 23063 7905 23075 7908
rect 23017 7899 23075 7905
rect 23658 7896 23664 7908
rect 23716 7896 23722 7948
rect 23768 7936 23796 7976
rect 26789 7973 26801 8007
rect 26835 8004 26847 8007
rect 27338 8004 27344 8016
rect 26835 7976 27344 8004
rect 26835 7973 26847 7976
rect 26789 7967 26847 7973
rect 27338 7964 27344 7976
rect 27396 7964 27402 8016
rect 27614 7964 27620 8016
rect 27672 8004 27678 8016
rect 27672 7976 29132 8004
rect 27672 7964 27678 7976
rect 27154 7936 27160 7948
rect 23768 7908 27160 7936
rect 27154 7896 27160 7908
rect 27212 7896 27218 7948
rect 27455 7939 27513 7945
rect 27455 7905 27467 7939
rect 27501 7936 27513 7939
rect 27706 7936 27712 7948
rect 27501 7908 27712 7936
rect 27501 7905 27513 7908
rect 27455 7899 27513 7905
rect 27706 7896 27712 7908
rect 27764 7896 27770 7948
rect 27798 7896 27804 7948
rect 27856 7936 27862 7948
rect 27856 7908 27901 7936
rect 27856 7896 27862 7908
rect 27982 7896 27988 7948
rect 28040 7936 28046 7948
rect 28994 7936 29000 7948
rect 28040 7908 28085 7936
rect 28955 7908 29000 7936
rect 28040 7896 28046 7908
rect 28994 7896 29000 7908
rect 29052 7896 29058 7948
rect 29104 7945 29132 7976
rect 29089 7939 29147 7945
rect 29089 7905 29101 7939
rect 29135 7905 29147 7939
rect 29089 7899 29147 7905
rect 19981 7871 20039 7877
rect 19981 7868 19993 7871
rect 19407 7840 19993 7868
rect 19981 7837 19993 7840
rect 20027 7868 20039 7871
rect 20530 7868 20536 7880
rect 20027 7840 20536 7868
rect 20027 7837 20039 7840
rect 19981 7831 20039 7837
rect 20530 7828 20536 7840
rect 20588 7828 20594 7880
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 21361 7871 21419 7877
rect 21361 7868 21373 7871
rect 20772 7840 21373 7868
rect 20772 7828 20778 7840
rect 21361 7837 21373 7840
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 22094 7828 22100 7880
rect 22152 7868 22158 7880
rect 22278 7868 22284 7880
rect 22152 7840 22284 7868
rect 22152 7828 22158 7840
rect 22278 7828 22284 7840
rect 22336 7828 22342 7880
rect 22922 7828 22928 7880
rect 22980 7868 22986 7880
rect 23109 7871 23167 7877
rect 23109 7868 23121 7871
rect 22980 7840 23121 7868
rect 22980 7828 22986 7840
rect 23109 7837 23121 7840
rect 23155 7837 23167 7871
rect 23109 7831 23167 7837
rect 27341 7871 27399 7877
rect 27341 7837 27353 7871
rect 27387 7868 27399 7871
rect 27387 7840 27660 7868
rect 27387 7837 27399 7840
rect 27341 7831 27399 7837
rect 2409 7803 2467 7809
rect 2409 7769 2421 7803
rect 2455 7800 2467 7803
rect 3142 7800 3148 7812
rect 2455 7772 3148 7800
rect 2455 7769 2467 7772
rect 2409 7763 2467 7769
rect 3142 7760 3148 7772
rect 3200 7760 3206 7812
rect 6638 7760 6644 7812
rect 6696 7800 6702 7812
rect 22462 7800 22468 7812
rect 6696 7772 22468 7800
rect 6696 7760 6702 7772
rect 22462 7760 22468 7772
rect 22520 7760 22526 7812
rect 22557 7803 22615 7809
rect 22557 7769 22569 7803
rect 22603 7800 22615 7803
rect 27632 7800 27660 7840
rect 27890 7828 27896 7880
rect 27948 7868 27954 7880
rect 27948 7840 30512 7868
rect 27948 7828 27954 7840
rect 30484 7809 30512 7840
rect 30469 7803 30527 7809
rect 22603 7772 24808 7800
rect 27632 7772 29316 7800
rect 22603 7769 22615 7772
rect 22557 7763 22615 7769
rect 11790 7732 11796 7744
rect 11751 7704 11796 7732
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 14274 7732 14280 7744
rect 14235 7704 14280 7732
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 15378 7692 15384 7744
rect 15436 7732 15442 7744
rect 15565 7735 15623 7741
rect 15565 7732 15577 7735
rect 15436 7704 15577 7732
rect 15436 7692 15442 7704
rect 15565 7701 15577 7704
rect 15611 7701 15623 7735
rect 15565 7695 15623 7701
rect 15654 7692 15660 7744
rect 15712 7732 15718 7744
rect 20346 7732 20352 7744
rect 15712 7704 20352 7732
rect 15712 7692 15718 7704
rect 20346 7692 20352 7704
rect 20404 7692 20410 7744
rect 24780 7732 24808 7772
rect 25682 7732 25688 7744
rect 24780 7704 25688 7732
rect 25682 7692 25688 7704
rect 25740 7692 25746 7744
rect 25774 7692 25780 7744
rect 25832 7732 25838 7744
rect 29288 7741 29316 7772
rect 30469 7769 30481 7803
rect 30515 7769 30527 7803
rect 30576 7800 30604 8044
rect 36004 8044 39712 8072
rect 31938 7964 31944 8016
rect 31996 8004 32002 8016
rect 33226 8004 33232 8016
rect 31996 7976 33232 8004
rect 31996 7964 32002 7976
rect 33226 7964 33232 7976
rect 33284 7964 33290 8016
rect 33410 7964 33416 8016
rect 33468 8004 33474 8016
rect 33873 8007 33931 8013
rect 33873 8004 33885 8007
rect 33468 7976 33885 8004
rect 33468 7964 33474 7976
rect 33873 7973 33885 7976
rect 33919 7973 33931 8007
rect 33873 7967 33931 7973
rect 30653 7939 30711 7945
rect 30653 7905 30665 7939
rect 30699 7905 30711 7939
rect 30653 7899 30711 7905
rect 31113 7939 31171 7945
rect 31113 7905 31125 7939
rect 31159 7936 31171 7939
rect 32030 7936 32036 7948
rect 31159 7908 32036 7936
rect 31159 7905 31171 7908
rect 31113 7899 31171 7905
rect 30668 7868 30696 7899
rect 32030 7896 32036 7908
rect 32088 7896 32094 7948
rect 32582 7936 32588 7948
rect 32543 7908 32588 7936
rect 32582 7896 32588 7908
rect 32640 7896 32646 7948
rect 34514 7936 34520 7948
rect 34475 7908 34520 7936
rect 34514 7896 34520 7908
rect 34572 7896 34578 7948
rect 34882 7936 34888 7948
rect 34843 7908 34888 7936
rect 34882 7896 34888 7908
rect 34940 7896 34946 7948
rect 34974 7896 34980 7948
rect 35032 7936 35038 7948
rect 36004 7945 36032 8044
rect 37366 7964 37372 8016
rect 37424 8004 37430 8016
rect 39574 8004 39580 8016
rect 37424 7976 39436 8004
rect 39535 7976 39580 8004
rect 37424 7964 37430 7976
rect 35989 7939 36047 7945
rect 35032 7908 35077 7936
rect 35032 7896 35038 7908
rect 35989 7905 36001 7939
rect 36035 7905 36047 7939
rect 35989 7899 36047 7905
rect 36078 7896 36084 7948
rect 36136 7936 36142 7948
rect 36262 7945 36268 7948
rect 36214 7939 36268 7945
rect 36136 7908 36181 7936
rect 36136 7896 36142 7908
rect 36214 7905 36226 7939
rect 36260 7905 36268 7939
rect 36214 7899 36268 7905
rect 36262 7896 36268 7899
rect 36320 7896 36326 7948
rect 37734 7936 37740 7948
rect 37695 7908 37740 7936
rect 37734 7896 37740 7908
rect 37792 7896 37798 7948
rect 39117 7939 39175 7945
rect 39117 7905 39129 7939
rect 39163 7936 39175 7939
rect 39298 7936 39304 7948
rect 39163 7908 39304 7936
rect 39163 7905 39175 7908
rect 39117 7899 39175 7905
rect 39298 7896 39304 7908
rect 39356 7896 39362 7948
rect 31386 7868 31392 7880
rect 30668 7840 31392 7868
rect 31386 7828 31392 7840
rect 31444 7828 31450 7880
rect 32398 7828 32404 7880
rect 32456 7868 32462 7880
rect 32493 7871 32551 7877
rect 32493 7868 32505 7871
rect 32456 7840 32505 7868
rect 32456 7828 32462 7840
rect 32493 7837 32505 7840
rect 32539 7868 32551 7871
rect 33778 7868 33784 7880
rect 32539 7840 33784 7868
rect 32539 7837 32551 7840
rect 32493 7831 32551 7837
rect 33778 7828 33784 7840
rect 33836 7828 33842 7880
rect 34425 7871 34483 7877
rect 34425 7837 34437 7871
rect 34471 7868 34483 7871
rect 36633 7871 36691 7877
rect 36633 7868 36645 7871
rect 34471 7840 36645 7868
rect 34471 7837 34483 7840
rect 34425 7831 34483 7837
rect 36633 7837 36645 7840
rect 36679 7837 36691 7871
rect 36633 7831 36691 7837
rect 38838 7828 38844 7880
rect 38896 7868 38902 7880
rect 39025 7871 39083 7877
rect 39025 7868 39037 7871
rect 38896 7840 39037 7868
rect 38896 7828 38902 7840
rect 39025 7837 39037 7840
rect 39071 7837 39083 7871
rect 39408 7868 39436 7976
rect 39574 7964 39580 7976
rect 39632 7964 39638 8016
rect 39684 8004 39712 8044
rect 39758 8032 39764 8084
rect 39816 8072 39822 8084
rect 39816 8044 44128 8072
rect 39816 8032 39822 8044
rect 42334 8004 42340 8016
rect 39684 7976 42340 8004
rect 42334 7964 42340 7976
rect 42392 7964 42398 8016
rect 43990 8004 43996 8016
rect 43640 7976 43996 8004
rect 40310 7896 40316 7948
rect 40368 7936 40374 7948
rect 40405 7939 40463 7945
rect 40405 7936 40417 7939
rect 40368 7908 40417 7936
rect 40368 7896 40374 7908
rect 40405 7905 40417 7908
rect 40451 7905 40463 7939
rect 40405 7899 40463 7905
rect 41141 7939 41199 7945
rect 41141 7905 41153 7939
rect 41187 7936 41199 7939
rect 41230 7936 41236 7948
rect 41187 7908 41236 7936
rect 41187 7905 41199 7908
rect 41141 7899 41199 7905
rect 41230 7896 41236 7908
rect 41288 7896 41294 7948
rect 41598 7896 41604 7948
rect 41656 7936 41662 7948
rect 41969 7939 42027 7945
rect 41969 7936 41981 7939
rect 41656 7908 41981 7936
rect 41656 7896 41662 7908
rect 41969 7905 41981 7908
rect 42015 7905 42027 7939
rect 41969 7899 42027 7905
rect 42242 7896 42248 7948
rect 42300 7936 42306 7948
rect 43530 7936 43536 7948
rect 42300 7908 43536 7936
rect 42300 7896 42306 7908
rect 43530 7896 43536 7908
rect 43588 7896 43594 7948
rect 43640 7945 43668 7976
rect 43990 7964 43996 7976
rect 44048 7964 44054 8016
rect 44100 7948 44128 8044
rect 44910 8032 44916 8084
rect 44968 8072 44974 8084
rect 46106 8072 46112 8084
rect 44968 8044 46112 8072
rect 44968 8032 44974 8044
rect 46106 8032 46112 8044
rect 46164 8032 46170 8084
rect 46198 8032 46204 8084
rect 46256 8072 46262 8084
rect 46477 8075 46535 8081
rect 46477 8072 46489 8075
rect 46256 8044 46489 8072
rect 46256 8032 46262 8044
rect 46477 8041 46489 8044
rect 46523 8041 46535 8075
rect 47762 8072 47768 8084
rect 47723 8044 47768 8072
rect 46477 8035 46535 8041
rect 47762 8032 47768 8044
rect 47820 8032 47826 8084
rect 55214 8072 55220 8084
rect 55175 8044 55220 8072
rect 55214 8032 55220 8044
rect 55272 8032 55278 8084
rect 56597 8075 56655 8081
rect 56597 8041 56609 8075
rect 56643 8072 56655 8075
rect 57238 8072 57244 8084
rect 56643 8044 57244 8072
rect 56643 8041 56655 8044
rect 56597 8035 56655 8041
rect 57238 8032 57244 8044
rect 57296 8032 57302 8084
rect 51718 8004 51724 8016
rect 46032 7976 51724 8004
rect 43625 7939 43683 7945
rect 43625 7905 43637 7939
rect 43671 7905 43683 7939
rect 44082 7936 44088 7948
rect 44043 7908 44088 7936
rect 43625 7899 43683 7905
rect 44082 7896 44088 7908
rect 44140 7896 44146 7948
rect 44450 7896 44456 7948
rect 44508 7936 44514 7948
rect 46032 7936 46060 7976
rect 51718 7964 51724 7976
rect 51776 7964 51782 8016
rect 55766 8004 55772 8016
rect 54772 7976 55772 8004
rect 44508 7908 46060 7936
rect 44508 7896 44514 7908
rect 46106 7896 46112 7948
rect 46164 7936 46170 7948
rect 47486 7936 47492 7948
rect 46164 7908 47492 7936
rect 46164 7896 46170 7908
rect 47486 7896 47492 7908
rect 47544 7936 47550 7948
rect 47581 7939 47639 7945
rect 47581 7936 47593 7939
rect 47544 7908 47593 7936
rect 47544 7896 47550 7908
rect 47581 7905 47593 7908
rect 47627 7905 47639 7939
rect 47581 7899 47639 7905
rect 50430 7896 50436 7948
rect 50488 7936 50494 7948
rect 51077 7939 51135 7945
rect 51077 7936 51089 7939
rect 50488 7908 51089 7936
rect 50488 7896 50494 7908
rect 51077 7905 51089 7908
rect 51123 7905 51135 7939
rect 51442 7936 51448 7948
rect 51403 7908 51448 7936
rect 51077 7899 51135 7905
rect 51442 7896 51448 7908
rect 51500 7896 51506 7948
rect 52454 7896 52460 7948
rect 52512 7936 52518 7948
rect 54772 7945 54800 7976
rect 55766 7964 55772 7976
rect 55824 7964 55830 8016
rect 58529 8007 58587 8013
rect 58529 7973 58541 8007
rect 58575 8004 58587 8007
rect 59262 8004 59268 8016
rect 58575 7976 59268 8004
rect 58575 7973 58587 7976
rect 58529 7967 58587 7973
rect 59262 7964 59268 7976
rect 59320 7964 59326 8016
rect 53193 7939 53251 7945
rect 53193 7936 53205 7939
rect 52512 7908 53205 7936
rect 52512 7896 52518 7908
rect 53193 7905 53205 7908
rect 53239 7905 53251 7939
rect 53193 7899 53251 7905
rect 54757 7939 54815 7945
rect 54757 7905 54769 7939
rect 54803 7905 54815 7939
rect 55030 7936 55036 7948
rect 54991 7908 55036 7936
rect 54757 7899 54815 7905
rect 55030 7896 55036 7908
rect 55088 7896 55094 7948
rect 55306 7896 55312 7948
rect 55364 7936 55370 7948
rect 56781 7939 56839 7945
rect 56781 7936 56793 7939
rect 55364 7908 56793 7936
rect 55364 7896 55370 7908
rect 56781 7905 56793 7908
rect 56827 7905 56839 7939
rect 56962 7936 56968 7948
rect 56923 7908 56968 7936
rect 56781 7899 56839 7905
rect 56962 7896 56968 7908
rect 57020 7896 57026 7948
rect 57333 7939 57391 7945
rect 57333 7936 57345 7939
rect 57072 7908 57345 7936
rect 44726 7868 44732 7880
rect 39408 7840 44732 7868
rect 39025 7831 39083 7837
rect 44726 7828 44732 7840
rect 44784 7828 44790 7880
rect 45005 7871 45063 7877
rect 45005 7837 45017 7871
rect 45051 7868 45063 7871
rect 45097 7871 45155 7877
rect 45097 7868 45109 7871
rect 45051 7840 45109 7868
rect 45051 7837 45063 7840
rect 45005 7831 45063 7837
rect 45097 7837 45109 7840
rect 45143 7868 45155 7871
rect 45278 7868 45284 7880
rect 45143 7840 45284 7868
rect 45143 7837 45155 7840
rect 45097 7831 45155 7837
rect 45278 7828 45284 7840
rect 45336 7828 45342 7880
rect 45373 7871 45431 7877
rect 45373 7837 45385 7871
rect 45419 7868 45431 7871
rect 45554 7868 45560 7880
rect 45419 7840 45560 7868
rect 45419 7837 45431 7840
rect 45373 7831 45431 7837
rect 45554 7828 45560 7840
rect 45612 7828 45618 7880
rect 45738 7828 45744 7880
rect 45796 7868 45802 7880
rect 49786 7868 49792 7880
rect 45796 7840 49792 7868
rect 45796 7828 45802 7840
rect 49786 7828 49792 7840
rect 49844 7828 49850 7880
rect 50798 7868 50804 7880
rect 50759 7840 50804 7868
rect 50798 7828 50804 7840
rect 50856 7828 50862 7880
rect 53098 7868 53104 7880
rect 53059 7840 53104 7868
rect 53098 7828 53104 7840
rect 53156 7828 53162 7880
rect 53653 7871 53711 7877
rect 53653 7837 53665 7871
rect 53699 7868 53711 7871
rect 55398 7868 55404 7880
rect 53699 7840 55404 7868
rect 53699 7837 53711 7840
rect 53653 7831 53711 7837
rect 55398 7828 55404 7840
rect 55456 7828 55462 7880
rect 55674 7828 55680 7880
rect 55732 7868 55738 7880
rect 57072 7868 57100 7908
rect 57333 7905 57345 7908
rect 57379 7905 57391 7939
rect 57333 7899 57391 7905
rect 58621 7939 58679 7945
rect 58621 7905 58633 7939
rect 58667 7905 58679 7939
rect 60274 7936 60280 7948
rect 60235 7908 60280 7936
rect 58621 7899 58679 7905
rect 57238 7868 57244 7880
rect 55732 7840 57100 7868
rect 57199 7840 57244 7868
rect 55732 7828 55738 7840
rect 57238 7828 57244 7840
rect 57296 7828 57302 7880
rect 57974 7828 57980 7880
rect 58032 7868 58038 7880
rect 58636 7868 58664 7899
rect 60274 7896 60280 7908
rect 60332 7896 60338 7948
rect 58032 7840 58664 7868
rect 58032 7828 58038 7840
rect 59446 7828 59452 7880
rect 59504 7868 59510 7880
rect 60185 7871 60243 7877
rect 60185 7868 60197 7871
rect 59504 7840 60197 7868
rect 59504 7828 59510 7840
rect 60185 7837 60197 7840
rect 60231 7837 60243 7871
rect 60185 7831 60243 7837
rect 30576 7772 32904 7800
rect 30469 7763 30527 7769
rect 28813 7735 28871 7741
rect 28813 7732 28825 7735
rect 25832 7704 28825 7732
rect 25832 7692 25838 7704
rect 28813 7701 28825 7704
rect 28859 7701 28871 7735
rect 28813 7695 28871 7701
rect 29273 7735 29331 7741
rect 29273 7701 29285 7735
rect 29319 7701 29331 7735
rect 29273 7695 29331 7701
rect 32306 7692 32312 7744
rect 32364 7732 32370 7744
rect 32769 7735 32827 7741
rect 32769 7732 32781 7735
rect 32364 7704 32781 7732
rect 32364 7692 32370 7704
rect 32769 7701 32781 7704
rect 32815 7701 32827 7735
rect 32876 7732 32904 7772
rect 33594 7760 33600 7812
rect 33652 7800 33658 7812
rect 42150 7800 42156 7812
rect 33652 7772 42012 7800
rect 42111 7772 42156 7800
rect 33652 7760 33658 7772
rect 37090 7732 37096 7744
rect 32876 7704 37096 7732
rect 32769 7695 32827 7701
rect 37090 7692 37096 7704
rect 37148 7692 37154 7744
rect 37921 7735 37979 7741
rect 37921 7701 37933 7735
rect 37967 7732 37979 7735
rect 38010 7732 38016 7744
rect 37967 7704 38016 7732
rect 37967 7701 37979 7704
rect 37921 7695 37979 7701
rect 38010 7692 38016 7704
rect 38068 7692 38074 7744
rect 40402 7692 40408 7744
rect 40460 7732 40466 7744
rect 40497 7735 40555 7741
rect 40497 7732 40509 7735
rect 40460 7704 40509 7732
rect 40460 7692 40466 7704
rect 40497 7701 40509 7704
rect 40543 7701 40555 7735
rect 41984 7732 42012 7772
rect 42150 7760 42156 7772
rect 42208 7760 42214 7812
rect 42260 7772 45140 7800
rect 42260 7732 42288 7772
rect 43438 7732 43444 7744
rect 41984 7704 42288 7732
rect 43399 7704 43444 7732
rect 40497 7695 40555 7701
rect 43438 7692 43444 7704
rect 43496 7692 43502 7744
rect 43530 7692 43536 7744
rect 43588 7732 43594 7744
rect 45005 7735 45063 7741
rect 45005 7732 45017 7735
rect 43588 7704 45017 7732
rect 43588 7692 43594 7704
rect 45005 7701 45017 7704
rect 45051 7701 45063 7735
rect 45112 7732 45140 7772
rect 51258 7760 51264 7812
rect 51316 7800 51322 7812
rect 51445 7803 51503 7809
rect 51445 7800 51457 7803
rect 51316 7772 51457 7800
rect 51316 7760 51322 7772
rect 51445 7769 51457 7772
rect 51491 7769 51503 7803
rect 53116 7800 53144 7828
rect 53742 7800 53748 7812
rect 53116 7772 53748 7800
rect 51445 7763 51503 7769
rect 53742 7760 53748 7772
rect 53800 7760 53806 7812
rect 54846 7800 54852 7812
rect 54807 7772 54852 7800
rect 54846 7760 54852 7772
rect 54904 7760 54910 7812
rect 47210 7732 47216 7744
rect 45112 7704 47216 7732
rect 45005 7695 45063 7701
rect 47210 7692 47216 7704
rect 47268 7692 47274 7744
rect 58342 7732 58348 7744
rect 58303 7704 58348 7732
rect 58342 7692 58348 7704
rect 58400 7692 58406 7744
rect 58802 7732 58808 7744
rect 58763 7704 58808 7732
rect 58802 7692 58808 7704
rect 58860 7692 58866 7744
rect 60458 7732 60464 7744
rect 60419 7704 60464 7732
rect 60458 7692 60464 7704
rect 60516 7692 60522 7744
rect 1104 7642 62192 7664
rect 1104 7590 11163 7642
rect 11215 7590 11227 7642
rect 11279 7590 11291 7642
rect 11343 7590 11355 7642
rect 11407 7590 31526 7642
rect 31578 7590 31590 7642
rect 31642 7590 31654 7642
rect 31706 7590 31718 7642
rect 31770 7590 51888 7642
rect 51940 7590 51952 7642
rect 52004 7590 52016 7642
rect 52068 7590 52080 7642
rect 52132 7590 62192 7642
rect 1104 7568 62192 7590
rect 5626 7528 5632 7540
rect 5587 7500 5632 7528
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 12713 7531 12771 7537
rect 12713 7497 12725 7531
rect 12759 7528 12771 7531
rect 13722 7528 13728 7540
rect 12759 7500 13728 7528
rect 12759 7497 12771 7500
rect 12713 7491 12771 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 14918 7488 14924 7540
rect 14976 7528 14982 7540
rect 16393 7531 16451 7537
rect 16393 7528 16405 7531
rect 14976 7500 16405 7528
rect 14976 7488 14982 7500
rect 16393 7497 16405 7500
rect 16439 7528 16451 7531
rect 16439 7500 19472 7528
rect 16439 7497 16451 7500
rect 16393 7491 16451 7497
rect 9766 7420 9772 7472
rect 9824 7460 9830 7472
rect 19444 7460 19472 7500
rect 19518 7488 19524 7540
rect 19576 7528 19582 7540
rect 19889 7531 19947 7537
rect 19889 7528 19901 7531
rect 19576 7500 19901 7528
rect 19576 7488 19582 7500
rect 19889 7497 19901 7500
rect 19935 7497 19947 7531
rect 19889 7491 19947 7497
rect 19978 7488 19984 7540
rect 20036 7528 20042 7540
rect 20036 7500 32444 7528
rect 20036 7488 20042 7500
rect 9824 7432 17264 7460
rect 19444 7432 20208 7460
rect 9824 7420 9830 7432
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7392 2927 7395
rect 3970 7392 3976 7404
rect 2915 7364 3976 7392
rect 2915 7361 2927 7364
rect 2869 7355 2927 7361
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 8110 7392 8116 7404
rect 5399 7364 8116 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7392 8355 7395
rect 8662 7392 8668 7404
rect 8343 7364 8668 7392
rect 8343 7361 8355 7364
rect 8297 7355 8355 7361
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 8754 7352 8760 7404
rect 8812 7392 8818 7404
rect 12986 7392 12992 7404
rect 8812 7364 10824 7392
rect 8812 7352 8818 7364
rect 3142 7324 3148 7336
rect 3103 7296 3148 7324
rect 3142 7284 3148 7296
rect 3200 7284 3206 7336
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7324 5503 7327
rect 6638 7324 6644 7336
rect 5491 7296 6644 7324
rect 5491 7293 5503 7296
rect 5445 7287 5503 7293
rect 4246 7216 4252 7268
rect 4304 7256 4310 7268
rect 5460 7256 5488 7287
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 8573 7327 8631 7333
rect 8573 7293 8585 7327
rect 8619 7324 8631 7327
rect 9674 7324 9680 7336
rect 8619 7296 9680 7324
rect 8619 7293 8631 7296
rect 8573 7287 8631 7293
rect 9674 7284 9680 7296
rect 9732 7284 9738 7336
rect 10796 7333 10824 7364
rect 11072 7364 12992 7392
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7293 10839 7327
rect 10781 7287 10839 7293
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 10962 7324 10968 7336
rect 10919 7296 10968 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11072 7333 11100 7364
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 15010 7392 15016 7404
rect 13648 7364 14872 7392
rect 14971 7364 15016 7392
rect 11057 7327 11115 7333
rect 11057 7293 11069 7327
rect 11103 7293 11115 7327
rect 12897 7327 12955 7333
rect 12897 7324 12909 7327
rect 11057 7287 11115 7293
rect 11900 7296 12909 7324
rect 9950 7256 9956 7268
rect 4304 7228 5488 7256
rect 9863 7228 9956 7256
rect 4304 7216 4310 7228
rect 9950 7216 9956 7228
rect 10008 7256 10014 7268
rect 11072 7256 11100 7287
rect 11900 7268 11928 7296
rect 12897 7293 12909 7296
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 13081 7327 13139 7333
rect 13081 7293 13093 7327
rect 13127 7324 13139 7327
rect 13354 7324 13360 7336
rect 13127 7296 13360 7324
rect 13127 7293 13139 7296
rect 13081 7287 13139 7293
rect 13354 7284 13360 7296
rect 13412 7284 13418 7336
rect 13446 7284 13452 7336
rect 13504 7324 13510 7336
rect 13648 7333 13676 7364
rect 13633 7327 13691 7333
rect 13504 7296 13549 7324
rect 13504 7284 13510 7296
rect 13633 7293 13645 7327
rect 13679 7293 13691 7327
rect 14458 7324 14464 7336
rect 14419 7296 14464 7324
rect 13633 7287 13691 7293
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 14642 7333 14648 7336
rect 14594 7327 14648 7333
rect 14594 7293 14606 7327
rect 14640 7293 14648 7327
rect 14594 7287 14648 7293
rect 14642 7284 14648 7287
rect 14700 7284 14706 7336
rect 14844 7324 14872 7364
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 16482 7392 16488 7404
rect 15856 7364 16488 7392
rect 15856 7324 15884 7364
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 17126 7392 17132 7404
rect 16592 7364 16896 7392
rect 17087 7364 17132 7392
rect 14844 7296 15884 7324
rect 15930 7284 15936 7336
rect 15988 7324 15994 7336
rect 16209 7327 16267 7333
rect 16209 7324 16221 7327
rect 15988 7296 16221 7324
rect 15988 7284 15994 7296
rect 16209 7293 16221 7296
rect 16255 7293 16267 7327
rect 16209 7287 16267 7293
rect 16301 7327 16359 7333
rect 16301 7293 16313 7327
rect 16347 7324 16359 7327
rect 16592 7324 16620 7364
rect 16758 7333 16764 7336
rect 16347 7296 16620 7324
rect 16710 7327 16764 7333
rect 16347 7293 16359 7296
rect 16301 7287 16359 7293
rect 16710 7293 16722 7327
rect 16756 7293 16764 7327
rect 16710 7287 16764 7293
rect 16758 7284 16764 7287
rect 16816 7284 16822 7336
rect 16868 7324 16896 7364
rect 17126 7352 17132 7364
rect 17184 7352 17190 7404
rect 17236 7392 17264 7432
rect 20070 7392 20076 7404
rect 17236 7364 20076 7392
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 16868 7296 18521 7324
rect 18509 7293 18521 7296
rect 18555 7293 18567 7327
rect 18782 7324 18788 7336
rect 18743 7296 18788 7324
rect 18509 7287 18567 7293
rect 18782 7284 18788 7296
rect 18840 7284 18846 7336
rect 10008 7228 11100 7256
rect 11517 7259 11575 7265
rect 10008 7216 10014 7228
rect 11517 7225 11529 7259
rect 11563 7256 11575 7259
rect 11882 7256 11888 7268
rect 11563 7228 11888 7256
rect 11563 7225 11575 7228
rect 11517 7219 11575 7225
rect 11882 7216 11888 7228
rect 11940 7216 11946 7268
rect 16577 7259 16635 7265
rect 16577 7225 16589 7259
rect 16623 7256 16635 7259
rect 17954 7256 17960 7268
rect 16623 7228 17960 7256
rect 16623 7225 16635 7228
rect 16577 7219 16635 7225
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 4430 7188 4436 7200
rect 4391 7160 4436 7188
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 13446 7148 13452 7200
rect 13504 7188 13510 7200
rect 15654 7188 15660 7200
rect 13504 7160 15660 7188
rect 13504 7148 13510 7160
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 16025 7191 16083 7197
rect 16025 7188 16037 7191
rect 15804 7160 16037 7188
rect 15804 7148 15810 7160
rect 16025 7157 16037 7160
rect 16071 7188 16083 7191
rect 16301 7191 16359 7197
rect 16301 7188 16313 7191
rect 16071 7160 16313 7188
rect 16071 7157 16083 7160
rect 16025 7151 16083 7157
rect 16301 7157 16313 7160
rect 16347 7157 16359 7191
rect 16301 7151 16359 7157
rect 16390 7148 16396 7200
rect 16448 7188 16454 7200
rect 19702 7188 19708 7200
rect 16448 7160 19708 7188
rect 16448 7148 16454 7160
rect 19702 7148 19708 7160
rect 19760 7148 19766 7200
rect 20180 7188 20208 7432
rect 20346 7420 20352 7472
rect 20404 7460 20410 7472
rect 20404 7432 22048 7460
rect 20404 7420 20410 7432
rect 20622 7352 20628 7404
rect 20680 7392 20686 7404
rect 20993 7395 21051 7401
rect 20993 7392 21005 7395
rect 20680 7364 21005 7392
rect 20680 7352 20686 7364
rect 20993 7361 21005 7364
rect 21039 7361 21051 7395
rect 20993 7355 21051 7361
rect 21545 7395 21603 7401
rect 21545 7361 21557 7395
rect 21591 7392 21603 7395
rect 21910 7392 21916 7404
rect 21591 7364 21916 7392
rect 21591 7361 21603 7364
rect 21545 7355 21603 7361
rect 21910 7352 21916 7364
rect 21968 7352 21974 7404
rect 22020 7392 22048 7432
rect 22278 7420 22284 7472
rect 22336 7460 22342 7472
rect 25774 7460 25780 7472
rect 22336 7432 25780 7460
rect 22336 7420 22342 7432
rect 25774 7420 25780 7432
rect 25832 7420 25838 7472
rect 27157 7463 27215 7469
rect 27157 7429 27169 7463
rect 27203 7460 27215 7463
rect 27982 7460 27988 7472
rect 27203 7432 27988 7460
rect 27203 7429 27215 7432
rect 27157 7423 27215 7429
rect 27982 7420 27988 7432
rect 28040 7420 28046 7472
rect 31386 7420 31392 7472
rect 31444 7460 31450 7472
rect 31938 7460 31944 7472
rect 31444 7432 31944 7460
rect 31444 7420 31450 7432
rect 31938 7420 31944 7432
rect 31996 7420 32002 7472
rect 32416 7460 32444 7500
rect 32490 7488 32496 7540
rect 32548 7528 32554 7540
rect 32548 7500 43484 7528
rect 32548 7488 32554 7500
rect 40310 7460 40316 7472
rect 32416 7432 40316 7460
rect 40310 7420 40316 7432
rect 40368 7420 40374 7472
rect 43456 7460 43484 7500
rect 44082 7488 44088 7540
rect 44140 7528 44146 7540
rect 44140 7500 55904 7528
rect 44140 7488 44146 7500
rect 47486 7460 47492 7472
rect 43456 7432 47072 7460
rect 32858 7392 32864 7404
rect 22020 7364 32864 7392
rect 21821 7327 21879 7333
rect 21821 7293 21833 7327
rect 21867 7293 21879 7327
rect 22002 7324 22008 7336
rect 21963 7296 22008 7324
rect 21821 7287 21879 7293
rect 20898 7216 20904 7268
rect 20956 7256 20962 7268
rect 21836 7256 21864 7287
rect 22002 7284 22008 7296
rect 22060 7284 22066 7336
rect 24210 7324 24216 7336
rect 24171 7296 24216 7324
rect 24210 7284 24216 7296
rect 24268 7284 24274 7336
rect 24305 7327 24363 7333
rect 24305 7293 24317 7327
rect 24351 7293 24363 7327
rect 24305 7287 24363 7293
rect 25593 7327 25651 7333
rect 25593 7293 25605 7327
rect 25639 7293 25651 7327
rect 25593 7287 25651 7293
rect 20956 7228 21864 7256
rect 20956 7216 20962 7228
rect 22462 7216 22468 7268
rect 22520 7256 22526 7268
rect 23290 7256 23296 7268
rect 22520 7228 23296 7256
rect 22520 7216 22526 7228
rect 23290 7216 23296 7228
rect 23348 7256 23354 7268
rect 24320 7256 24348 7287
rect 23348 7228 24348 7256
rect 24765 7259 24823 7265
rect 23348 7216 23354 7228
rect 24765 7225 24777 7259
rect 24811 7256 24823 7259
rect 25038 7256 25044 7268
rect 24811 7228 25044 7256
rect 24811 7225 24823 7228
rect 24765 7219 24823 7225
rect 25038 7216 25044 7228
rect 25096 7216 25102 7268
rect 25608 7200 25636 7287
rect 27154 7284 27160 7336
rect 27212 7324 27218 7336
rect 27341 7327 27399 7333
rect 27341 7324 27353 7327
rect 27212 7296 27353 7324
rect 27212 7284 27218 7296
rect 27341 7293 27353 7296
rect 27387 7293 27399 7327
rect 27341 7287 27399 7293
rect 27430 7284 27436 7336
rect 27488 7324 27494 7336
rect 27709 7327 27767 7333
rect 27709 7324 27721 7327
rect 27488 7296 27721 7324
rect 27488 7284 27494 7296
rect 27709 7293 27721 7296
rect 27755 7293 27767 7327
rect 27709 7287 27767 7293
rect 27801 7327 27859 7333
rect 27801 7293 27813 7327
rect 27847 7324 27859 7327
rect 28994 7324 29000 7336
rect 27847 7296 29000 7324
rect 27847 7293 27859 7296
rect 27801 7287 27859 7293
rect 28994 7284 29000 7296
rect 29052 7284 29058 7336
rect 29457 7327 29515 7333
rect 29457 7293 29469 7327
rect 29503 7324 29515 7327
rect 29546 7324 29552 7336
rect 29503 7296 29552 7324
rect 29503 7293 29515 7296
rect 29457 7287 29515 7293
rect 29546 7284 29552 7296
rect 29604 7284 29610 7336
rect 30668 7333 30696 7364
rect 32858 7352 32864 7364
rect 32916 7352 32922 7404
rect 33594 7392 33600 7404
rect 33555 7364 33600 7392
rect 33594 7352 33600 7364
rect 33652 7352 33658 7404
rect 33778 7352 33784 7404
rect 33836 7392 33842 7404
rect 36354 7392 36360 7404
rect 33836 7364 36360 7392
rect 33836 7352 33842 7364
rect 36354 7352 36360 7364
rect 36412 7392 36418 7404
rect 36412 7364 36676 7392
rect 36412 7352 36418 7364
rect 30653 7327 30711 7333
rect 30653 7293 30665 7327
rect 30699 7293 30711 7327
rect 30653 7287 30711 7293
rect 31757 7327 31815 7333
rect 31757 7293 31769 7327
rect 31803 7324 31815 7327
rect 32582 7324 32588 7336
rect 31803 7296 32588 7324
rect 31803 7293 31815 7296
rect 31757 7287 31815 7293
rect 32582 7284 32588 7296
rect 32640 7284 32646 7336
rect 33226 7324 33232 7336
rect 33187 7296 33232 7324
rect 33226 7284 33232 7296
rect 33284 7284 33290 7336
rect 33965 7327 34023 7333
rect 33965 7293 33977 7327
rect 34011 7324 34023 7327
rect 34330 7324 34336 7336
rect 34011 7296 34336 7324
rect 34011 7293 34023 7296
rect 33965 7287 34023 7293
rect 34330 7284 34336 7296
rect 34388 7284 34394 7336
rect 35526 7324 35532 7336
rect 35487 7296 35532 7324
rect 35526 7284 35532 7296
rect 35584 7284 35590 7336
rect 36078 7324 36084 7336
rect 36039 7296 36084 7324
rect 36078 7284 36084 7296
rect 36136 7284 36142 7336
rect 36170 7284 36176 7336
rect 36228 7324 36234 7336
rect 36648 7333 36676 7364
rect 38102 7352 38108 7404
rect 38160 7392 38166 7404
rect 38562 7392 38568 7404
rect 38160 7364 38568 7392
rect 38160 7352 38166 7364
rect 38562 7352 38568 7364
rect 38620 7352 38626 7404
rect 40678 7392 40684 7404
rect 39224 7364 40684 7392
rect 36265 7327 36323 7333
rect 36265 7324 36277 7327
rect 36228 7296 36277 7324
rect 36228 7284 36234 7296
rect 36265 7293 36277 7296
rect 36311 7293 36323 7327
rect 36265 7287 36323 7293
rect 36633 7327 36691 7333
rect 36633 7293 36645 7327
rect 36679 7293 36691 7327
rect 36998 7324 37004 7336
rect 36959 7296 37004 7324
rect 36633 7287 36691 7293
rect 36998 7284 37004 7296
rect 37056 7284 37062 7336
rect 37090 7284 37096 7336
rect 37148 7324 37154 7336
rect 39224 7333 39252 7364
rect 40678 7352 40684 7364
rect 40736 7352 40742 7404
rect 41325 7395 41383 7401
rect 41325 7361 41337 7395
rect 41371 7392 41383 7395
rect 42886 7392 42892 7404
rect 41371 7364 42892 7392
rect 41371 7361 41383 7364
rect 41325 7355 41383 7361
rect 42886 7352 42892 7364
rect 42944 7352 42950 7404
rect 44177 7395 44235 7401
rect 44177 7361 44189 7395
rect 44223 7392 44235 7395
rect 44266 7392 44272 7404
rect 44223 7364 44272 7392
rect 44223 7361 44235 7364
rect 44177 7355 44235 7361
rect 44266 7352 44272 7364
rect 44324 7352 44330 7404
rect 44726 7392 44732 7404
rect 44687 7364 44732 7392
rect 44726 7352 44732 7364
rect 44784 7352 44790 7404
rect 46382 7392 46388 7404
rect 45020 7364 46388 7392
rect 39209 7327 39267 7333
rect 39209 7324 39221 7327
rect 37148 7296 39221 7324
rect 37148 7284 37154 7296
rect 39209 7293 39221 7296
rect 39255 7293 39267 7327
rect 39209 7287 39267 7293
rect 39577 7327 39635 7333
rect 39577 7293 39589 7327
rect 39623 7324 39635 7327
rect 41233 7327 41291 7333
rect 41233 7324 41245 7327
rect 39623 7296 41245 7324
rect 39623 7293 39635 7296
rect 39577 7287 39635 7293
rect 41233 7293 41245 7296
rect 41279 7293 41291 7327
rect 42061 7327 42119 7333
rect 42061 7324 42073 7327
rect 41233 7287 41291 7293
rect 41340 7296 42073 7324
rect 41340 7268 41368 7296
rect 42061 7293 42073 7296
rect 42107 7293 42119 7327
rect 42061 7287 42119 7293
rect 42150 7284 42156 7336
rect 42208 7324 42214 7336
rect 43070 7324 43076 7336
rect 42208 7296 42253 7324
rect 43031 7296 43076 7324
rect 42208 7284 42214 7296
rect 43070 7284 43076 7296
rect 43128 7284 43134 7336
rect 43990 7284 43996 7336
rect 44048 7324 44054 7336
rect 45020 7333 45048 7364
rect 46382 7352 46388 7364
rect 46440 7352 46446 7404
rect 45005 7327 45063 7333
rect 45005 7324 45017 7327
rect 44048 7296 45017 7324
rect 44048 7284 44054 7296
rect 45005 7293 45017 7296
rect 45051 7293 45063 7327
rect 45186 7324 45192 7336
rect 45147 7296 45192 7324
rect 45005 7287 45063 7293
rect 45186 7284 45192 7296
rect 45244 7284 45250 7336
rect 46198 7284 46204 7336
rect 46256 7324 46262 7336
rect 46661 7327 46719 7333
rect 46661 7324 46673 7327
rect 46256 7296 46673 7324
rect 46256 7284 46262 7296
rect 46661 7293 46673 7296
rect 46707 7293 46719 7327
rect 46661 7287 46719 7293
rect 46937 7327 46995 7333
rect 46937 7293 46949 7327
rect 46983 7293 46995 7327
rect 47044 7324 47072 7432
rect 47136 7432 47492 7460
rect 47136 7401 47164 7432
rect 47486 7420 47492 7432
rect 47544 7420 47550 7472
rect 47121 7395 47179 7401
rect 47121 7361 47133 7395
rect 47167 7361 47179 7395
rect 47121 7355 47179 7361
rect 47210 7352 47216 7404
rect 47268 7392 47274 7404
rect 54754 7392 54760 7404
rect 47268 7364 54760 7392
rect 47268 7352 47274 7364
rect 54754 7352 54760 7364
rect 54812 7352 54818 7404
rect 55876 7336 55904 7500
rect 56045 7395 56103 7401
rect 56045 7361 56057 7395
rect 56091 7392 56103 7395
rect 56962 7392 56968 7404
rect 56091 7364 56968 7392
rect 56091 7361 56103 7364
rect 56045 7355 56103 7361
rect 56962 7352 56968 7364
rect 57020 7352 57026 7404
rect 58066 7352 58072 7404
rect 58124 7392 58130 7404
rect 58434 7392 58440 7404
rect 58124 7364 58440 7392
rect 58124 7352 58130 7364
rect 58434 7352 58440 7364
rect 58492 7392 58498 7404
rect 58529 7395 58587 7401
rect 58529 7392 58541 7395
rect 58492 7364 58541 7392
rect 58492 7352 58498 7364
rect 58529 7361 58541 7364
rect 58575 7361 58587 7395
rect 58529 7355 58587 7361
rect 48685 7327 48743 7333
rect 48685 7324 48697 7327
rect 47044 7296 48697 7324
rect 46937 7287 46995 7293
rect 48685 7293 48697 7296
rect 48731 7324 48743 7327
rect 50525 7327 50583 7333
rect 50525 7324 50537 7327
rect 48731 7296 50537 7324
rect 48731 7293 48743 7296
rect 48685 7287 48743 7293
rect 50525 7293 50537 7296
rect 50571 7293 50583 7327
rect 50525 7287 50583 7293
rect 29273 7259 29331 7265
rect 29273 7225 29285 7259
rect 29319 7256 29331 7259
rect 33042 7256 33048 7268
rect 29319 7228 33048 7256
rect 29319 7225 29331 7228
rect 29273 7219 29331 7225
rect 33042 7216 33048 7228
rect 33100 7216 33106 7268
rect 35342 7216 35348 7268
rect 35400 7256 35406 7268
rect 35713 7259 35771 7265
rect 35713 7256 35725 7259
rect 35400 7228 35725 7256
rect 35400 7216 35406 7228
rect 35713 7225 35725 7228
rect 35759 7256 35771 7259
rect 37274 7256 37280 7268
rect 35759 7228 37280 7256
rect 35759 7225 35771 7228
rect 35713 7219 35771 7225
rect 37274 7216 37280 7228
rect 37332 7216 37338 7268
rect 38746 7216 38752 7268
rect 38804 7256 38810 7268
rect 39022 7259 39080 7265
rect 39022 7256 39034 7259
rect 38804 7228 39034 7256
rect 38804 7216 38810 7228
rect 39022 7225 39034 7228
rect 39068 7256 39080 7259
rect 39068 7228 39896 7256
rect 39068 7225 39080 7228
rect 39022 7219 39080 7225
rect 25590 7188 25596 7200
rect 20180 7160 25596 7188
rect 25590 7148 25596 7160
rect 25648 7148 25654 7200
rect 28994 7148 29000 7200
rect 29052 7188 29058 7200
rect 29549 7191 29607 7197
rect 29549 7188 29561 7191
rect 29052 7160 29561 7188
rect 29052 7148 29058 7160
rect 29549 7157 29561 7160
rect 29595 7157 29607 7191
rect 29549 7151 29607 7157
rect 30466 7148 30472 7200
rect 30524 7188 30530 7200
rect 30834 7188 30840 7200
rect 30524 7160 30840 7188
rect 30524 7148 30530 7160
rect 30834 7148 30840 7160
rect 30892 7148 30898 7200
rect 33778 7148 33784 7200
rect 33836 7188 33842 7200
rect 35434 7188 35440 7200
rect 33836 7160 35440 7188
rect 33836 7148 33842 7160
rect 35434 7148 35440 7160
rect 35492 7188 35498 7200
rect 38562 7188 38568 7200
rect 35492 7160 38568 7188
rect 35492 7148 35498 7160
rect 38562 7148 38568 7160
rect 38620 7148 38626 7200
rect 39868 7188 39896 7228
rect 41322 7216 41328 7268
rect 41380 7216 41386 7268
rect 43346 7256 43352 7268
rect 41432 7228 43352 7256
rect 41432 7188 41460 7228
rect 43346 7216 43352 7228
rect 43404 7216 43410 7268
rect 46106 7256 46112 7268
rect 46067 7228 46112 7256
rect 46106 7216 46112 7228
rect 46164 7216 46170 7268
rect 46952 7256 46980 7287
rect 51534 7284 51540 7336
rect 51592 7324 51598 7336
rect 51718 7324 51724 7336
rect 51592 7296 51724 7324
rect 51592 7284 51598 7296
rect 51718 7284 51724 7296
rect 51776 7324 51782 7336
rect 52273 7327 52331 7333
rect 52273 7324 52285 7327
rect 51776 7296 52285 7324
rect 51776 7284 51782 7296
rect 52273 7293 52285 7296
rect 52319 7293 52331 7327
rect 52546 7324 52552 7336
rect 52507 7296 52552 7324
rect 52273 7287 52331 7293
rect 52546 7284 52552 7296
rect 52604 7284 52610 7336
rect 55766 7324 55772 7336
rect 55727 7296 55772 7324
rect 55766 7284 55772 7296
rect 55824 7284 55830 7336
rect 55858 7284 55864 7336
rect 55916 7324 55922 7336
rect 56229 7327 56287 7333
rect 56229 7324 56241 7327
rect 55916 7296 56241 7324
rect 55916 7284 55922 7296
rect 56229 7293 56241 7296
rect 56275 7293 56287 7327
rect 56229 7287 56287 7293
rect 57333 7327 57391 7333
rect 57333 7293 57345 7327
rect 57379 7293 57391 7327
rect 57333 7287 57391 7293
rect 50430 7256 50436 7268
rect 46952 7228 50436 7256
rect 50430 7216 50436 7228
rect 50488 7216 50494 7268
rect 53926 7256 53932 7268
rect 53887 7228 53932 7256
rect 53926 7216 53932 7228
rect 53984 7216 53990 7268
rect 54754 7216 54760 7268
rect 54812 7256 54818 7268
rect 57348 7256 57376 7287
rect 58618 7284 58624 7336
rect 58676 7324 58682 7336
rect 58805 7327 58863 7333
rect 58805 7324 58817 7327
rect 58676 7296 58817 7324
rect 58676 7284 58682 7296
rect 58805 7293 58817 7296
rect 58851 7293 58863 7327
rect 58805 7287 58863 7293
rect 54812 7228 57376 7256
rect 54812 7216 54818 7228
rect 39868 7160 41460 7188
rect 42150 7148 42156 7200
rect 42208 7188 42214 7200
rect 43257 7191 43315 7197
rect 43257 7188 43269 7191
rect 42208 7160 43269 7188
rect 42208 7148 42214 7160
rect 43257 7157 43269 7160
rect 43303 7157 43315 7191
rect 43257 7151 43315 7157
rect 44726 7148 44732 7200
rect 44784 7188 44790 7200
rect 47210 7188 47216 7200
rect 44784 7160 47216 7188
rect 44784 7148 44790 7160
rect 47210 7148 47216 7160
rect 47268 7148 47274 7200
rect 48222 7148 48228 7200
rect 48280 7188 48286 7200
rect 48869 7191 48927 7197
rect 48869 7188 48881 7191
rect 48280 7160 48881 7188
rect 48280 7148 48286 7160
rect 48869 7157 48881 7160
rect 48915 7157 48927 7191
rect 48869 7151 48927 7157
rect 50709 7191 50767 7197
rect 50709 7157 50721 7191
rect 50755 7188 50767 7191
rect 53190 7188 53196 7200
rect 50755 7160 53196 7188
rect 50755 7157 50767 7160
rect 50709 7151 50767 7157
rect 53190 7148 53196 7160
rect 53248 7148 53254 7200
rect 56962 7148 56968 7200
rect 57020 7188 57026 7200
rect 57517 7191 57575 7197
rect 57517 7188 57529 7191
rect 57020 7160 57529 7188
rect 57020 7148 57026 7160
rect 57517 7157 57529 7160
rect 57563 7157 57575 7191
rect 59906 7188 59912 7200
rect 59867 7160 59912 7188
rect 57517 7151 57575 7157
rect 59906 7148 59912 7160
rect 59964 7148 59970 7200
rect 1104 7098 62192 7120
rect 1104 7046 21344 7098
rect 21396 7046 21408 7098
rect 21460 7046 21472 7098
rect 21524 7046 21536 7098
rect 21588 7046 41707 7098
rect 41759 7046 41771 7098
rect 41823 7046 41835 7098
rect 41887 7046 41899 7098
rect 41951 7046 62192 7098
rect 1104 7024 62192 7046
rect 3050 6984 3056 6996
rect 3011 6956 3056 6984
rect 3050 6944 3056 6956
rect 3108 6944 3114 6996
rect 34241 6987 34299 6993
rect 34241 6984 34253 6987
rect 4172 6956 34253 6984
rect 4172 6916 4200 6956
rect 34241 6953 34253 6956
rect 34287 6953 34299 6987
rect 37182 6984 37188 6996
rect 34241 6947 34299 6953
rect 34348 6956 37188 6984
rect 8754 6916 8760 6928
rect 2976 6888 4200 6916
rect 8496 6888 8760 6916
rect 2976 6857 3004 6888
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6817 3019 6851
rect 2961 6811 3019 6817
rect 3970 6808 3976 6860
rect 4028 6848 4034 6860
rect 4065 6851 4123 6857
rect 4065 6848 4077 6851
rect 4028 6820 4077 6848
rect 4028 6808 4034 6820
rect 4065 6817 4077 6820
rect 4111 6848 4123 6851
rect 4154 6848 4160 6860
rect 4111 6820 4160 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 4154 6808 4160 6820
rect 4212 6808 4218 6860
rect 5718 6848 5724 6860
rect 5631 6820 5724 6848
rect 5718 6808 5724 6820
rect 5776 6848 5782 6860
rect 6454 6848 6460 6860
rect 5776 6820 6460 6848
rect 5776 6808 5782 6820
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 6638 6848 6644 6860
rect 6599 6820 6644 6848
rect 6638 6808 6644 6820
rect 6696 6808 6702 6860
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6848 8263 6851
rect 8496 6848 8524 6888
rect 8754 6876 8760 6888
rect 8812 6876 8818 6928
rect 10042 6916 10048 6928
rect 9600 6888 10048 6916
rect 8251 6820 8524 6848
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 8570 6808 8576 6860
rect 8628 6848 8634 6860
rect 9600 6848 9628 6888
rect 10042 6876 10048 6888
rect 10100 6876 10106 6928
rect 16114 6916 16120 6928
rect 10612 6888 16120 6916
rect 10612 6860 10640 6888
rect 16114 6876 16120 6888
rect 16172 6876 16178 6928
rect 17681 6919 17739 6925
rect 17681 6885 17693 6919
rect 17727 6916 17739 6919
rect 18046 6916 18052 6928
rect 17727 6888 18052 6916
rect 17727 6885 17739 6888
rect 17681 6879 17739 6885
rect 18046 6876 18052 6888
rect 18104 6876 18110 6928
rect 18693 6919 18751 6925
rect 18693 6885 18705 6919
rect 18739 6916 18751 6919
rect 18782 6916 18788 6928
rect 18739 6888 18788 6916
rect 18739 6885 18751 6888
rect 18693 6879 18751 6885
rect 18782 6876 18788 6888
rect 18840 6876 18846 6928
rect 20254 6916 20260 6928
rect 19352 6888 20260 6916
rect 8628 6820 9628 6848
rect 9677 6851 9735 6857
rect 8628 6808 8634 6820
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 9950 6848 9956 6860
rect 9723 6820 9956 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 10594 6848 10600 6860
rect 10507 6820 10600 6848
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 11882 6848 11888 6860
rect 11843 6820 11888 6848
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 12158 6808 12164 6860
rect 12216 6848 12222 6860
rect 12575 6851 12633 6857
rect 12575 6848 12587 6851
rect 12216 6820 12587 6848
rect 12216 6808 12222 6820
rect 12575 6817 12587 6820
rect 12621 6817 12633 6851
rect 12575 6811 12633 6817
rect 12713 6851 12771 6857
rect 12713 6817 12725 6851
rect 12759 6817 12771 6851
rect 13814 6848 13820 6860
rect 13775 6820 13820 6848
rect 12713 6811 12771 6817
rect 4338 6780 4344 6792
rect 4299 6752 4344 6780
rect 4338 6740 4344 6752
rect 4396 6740 4402 6792
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6780 6607 6783
rect 7742 6780 7748 6792
rect 6595 6752 7748 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6780 8447 6783
rect 10318 6780 10324 6792
rect 8435 6752 10324 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 10318 6740 10324 6752
rect 10376 6780 10382 6792
rect 10689 6783 10747 6789
rect 10689 6780 10701 6783
rect 10376 6752 10701 6780
rect 10376 6740 10382 6752
rect 10689 6749 10701 6752
rect 10735 6749 10747 6783
rect 10689 6743 10747 6749
rect 11974 6740 11980 6792
rect 12032 6780 12038 6792
rect 12032 6752 12077 6780
rect 12032 6740 12038 6752
rect 10134 6712 10140 6724
rect 10095 6684 10140 6712
rect 10134 6672 10140 6684
rect 10192 6672 10198 6724
rect 12728 6712 12756 6811
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 14001 6851 14059 6857
rect 14001 6817 14013 6851
rect 14047 6848 14059 6851
rect 14090 6848 14096 6860
rect 14047 6820 14096 6848
rect 14047 6817 14059 6820
rect 14001 6811 14059 6817
rect 14090 6808 14096 6820
rect 14148 6848 14154 6860
rect 15102 6848 15108 6860
rect 14148 6820 15108 6848
rect 14148 6808 14154 6820
rect 15102 6808 15108 6820
rect 15160 6808 15166 6860
rect 19352 6857 19380 6888
rect 20254 6876 20260 6888
rect 20312 6876 20318 6928
rect 24872 6888 25176 6916
rect 19337 6851 19395 6857
rect 19337 6848 19349 6851
rect 15212 6820 19349 6848
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 15212 6780 15240 6820
rect 19337 6817 19349 6820
rect 19383 6817 19395 6851
rect 19702 6848 19708 6860
rect 19663 6820 19708 6848
rect 19337 6811 19395 6817
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 20898 6848 20904 6860
rect 20859 6820 20904 6848
rect 20898 6808 20904 6820
rect 20956 6808 20962 6860
rect 20990 6808 20996 6860
rect 21048 6848 21054 6860
rect 21453 6851 21511 6857
rect 21453 6848 21465 6851
rect 21048 6820 21465 6848
rect 21048 6808 21054 6820
rect 21453 6817 21465 6820
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 22925 6851 22983 6857
rect 22925 6817 22937 6851
rect 22971 6817 22983 6851
rect 23382 6848 23388 6860
rect 23343 6820 23388 6848
rect 22925 6811 22983 6817
rect 13136 6752 15240 6780
rect 13136 6740 13142 6752
rect 15746 6740 15752 6792
rect 15804 6780 15810 6792
rect 16025 6783 16083 6789
rect 16025 6780 16037 6783
rect 15804 6752 16037 6780
rect 15804 6740 15810 6752
rect 16025 6749 16037 6752
rect 16071 6749 16083 6783
rect 16298 6780 16304 6792
rect 16259 6752 16304 6780
rect 16025 6743 16083 6749
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 19242 6780 19248 6792
rect 19203 6752 19248 6780
rect 19242 6740 19248 6752
rect 19300 6740 19306 6792
rect 19518 6740 19524 6792
rect 19576 6780 19582 6792
rect 19797 6783 19855 6789
rect 19797 6780 19809 6783
rect 19576 6752 19809 6780
rect 19576 6740 19582 6752
rect 19797 6749 19809 6752
rect 19843 6749 19855 6783
rect 19797 6743 19855 6749
rect 22370 6740 22376 6792
rect 22428 6780 22434 6792
rect 22833 6783 22891 6789
rect 22833 6780 22845 6783
rect 22428 6752 22845 6780
rect 22428 6740 22434 6752
rect 22833 6749 22845 6752
rect 22879 6749 22891 6783
rect 22940 6780 22968 6811
rect 23382 6808 23388 6820
rect 23440 6808 23446 6860
rect 23566 6808 23572 6860
rect 23624 6848 23630 6860
rect 24872 6848 24900 6888
rect 25038 6848 25044 6860
rect 23624 6820 24900 6848
rect 24999 6820 25044 6848
rect 23624 6808 23630 6820
rect 25038 6808 25044 6820
rect 25096 6808 25102 6860
rect 25148 6848 25176 6888
rect 25332 6888 25544 6916
rect 25225 6851 25283 6857
rect 25225 6848 25237 6851
rect 25148 6820 25237 6848
rect 25225 6817 25237 6820
rect 25271 6848 25283 6851
rect 25332 6848 25360 6888
rect 25271 6820 25360 6848
rect 25409 6851 25467 6857
rect 25271 6817 25283 6820
rect 25225 6811 25283 6817
rect 25409 6817 25421 6851
rect 25455 6817 25467 6851
rect 25516 6848 25544 6888
rect 25682 6876 25688 6928
rect 25740 6916 25746 6928
rect 27154 6916 27160 6928
rect 25740 6888 27016 6916
rect 27115 6888 27160 6916
rect 25740 6876 25746 6888
rect 26988 6860 27016 6888
rect 27154 6876 27160 6888
rect 27212 6876 27218 6928
rect 34348 6916 34376 6956
rect 37182 6944 37188 6956
rect 37240 6944 37246 6996
rect 37734 6944 37740 6996
rect 37792 6984 37798 6996
rect 37829 6987 37887 6993
rect 37829 6984 37841 6987
rect 37792 6956 37841 6984
rect 37792 6944 37798 6956
rect 37829 6953 37841 6956
rect 37875 6953 37887 6987
rect 37829 6947 37887 6953
rect 45554 6944 45560 6996
rect 45612 6984 45618 6996
rect 45649 6987 45707 6993
rect 45649 6984 45661 6987
rect 45612 6956 45661 6984
rect 45612 6944 45618 6956
rect 45649 6953 45661 6956
rect 45695 6953 45707 6987
rect 45649 6947 45707 6953
rect 51000 6956 56824 6984
rect 29748 6888 29960 6916
rect 26878 6848 26884 6860
rect 25516 6820 26884 6848
rect 25409 6811 25467 6817
rect 23842 6780 23848 6792
rect 22940 6752 23848 6780
rect 22833 6743 22891 6749
rect 23842 6740 23848 6752
rect 23900 6740 23906 6792
rect 25424 6780 25452 6811
rect 26878 6808 26884 6820
rect 26936 6808 26942 6860
rect 26970 6808 26976 6860
rect 27028 6848 27034 6860
rect 27525 6851 27583 6857
rect 27028 6820 27121 6848
rect 27028 6808 27034 6820
rect 27525 6817 27537 6851
rect 27571 6848 27583 6851
rect 27798 6848 27804 6860
rect 27571 6820 27804 6848
rect 27571 6817 27583 6820
rect 27525 6811 27583 6817
rect 27798 6808 27804 6820
rect 27856 6808 27862 6860
rect 27982 6848 27988 6860
rect 27943 6820 27988 6848
rect 27982 6808 27988 6820
rect 28040 6808 28046 6860
rect 28074 6808 28080 6860
rect 28132 6848 28138 6860
rect 28132 6820 28225 6848
rect 28132 6808 28138 6820
rect 28258 6808 28264 6860
rect 28316 6848 28322 6860
rect 28445 6851 28503 6857
rect 28445 6848 28457 6851
rect 28316 6820 28457 6848
rect 28316 6808 28322 6820
rect 28445 6817 28457 6820
rect 28491 6817 28503 6851
rect 28445 6811 28503 6817
rect 25958 6780 25964 6792
rect 25424 6752 25964 6780
rect 25958 6740 25964 6752
rect 26016 6740 26022 6792
rect 14458 6712 14464 6724
rect 12728 6684 14464 6712
rect 14458 6672 14464 6684
rect 14516 6672 14522 6724
rect 17954 6672 17960 6724
rect 18012 6712 18018 6724
rect 20993 6715 21051 6721
rect 20993 6712 21005 6715
rect 18012 6684 21005 6712
rect 18012 6672 18018 6684
rect 20993 6681 21005 6684
rect 21039 6681 21051 6715
rect 20993 6675 21051 6681
rect 24857 6715 24915 6721
rect 24857 6681 24869 6715
rect 24903 6712 24915 6715
rect 25222 6712 25228 6724
rect 24903 6684 25228 6712
rect 24903 6681 24915 6684
rect 24857 6675 24915 6681
rect 25222 6672 25228 6684
rect 25280 6672 25286 6724
rect 27522 6672 27528 6724
rect 27580 6712 27586 6724
rect 28092 6712 28120 6808
rect 28460 6780 28488 6811
rect 28534 6808 28540 6860
rect 28592 6848 28598 6860
rect 29748 6848 29776 6888
rect 28592 6820 29776 6848
rect 29825 6851 29883 6857
rect 28592 6808 28598 6820
rect 29825 6817 29837 6851
rect 29871 6817 29883 6851
rect 29932 6848 29960 6888
rect 33704 6888 34376 6916
rect 30558 6848 30564 6860
rect 29932 6820 30564 6848
rect 29825 6811 29883 6817
rect 28718 6780 28724 6792
rect 28460 6752 28724 6780
rect 28718 6740 28724 6752
rect 28776 6740 28782 6792
rect 29840 6780 29868 6811
rect 30558 6808 30564 6820
rect 30616 6808 30622 6860
rect 30650 6808 30656 6860
rect 30708 6848 30714 6860
rect 30929 6851 30987 6857
rect 30929 6848 30941 6851
rect 30708 6820 30941 6848
rect 30708 6808 30714 6820
rect 30929 6817 30941 6820
rect 30975 6848 30987 6851
rect 32306 6848 32312 6860
rect 30975 6820 32312 6848
rect 30975 6817 30987 6820
rect 30929 6811 30987 6817
rect 32306 6808 32312 6820
rect 32364 6808 32370 6860
rect 32674 6848 32680 6860
rect 32635 6820 32680 6848
rect 32674 6808 32680 6820
rect 32732 6848 32738 6860
rect 33410 6848 33416 6860
rect 32732 6820 33416 6848
rect 32732 6808 32738 6820
rect 33410 6808 33416 6820
rect 33468 6808 33474 6860
rect 32692 6780 32720 6808
rect 33704 6780 33732 6888
rect 41230 6876 41236 6928
rect 41288 6916 41294 6928
rect 51000 6916 51028 6956
rect 51350 6916 51356 6928
rect 41288 6888 51028 6916
rect 51092 6888 51356 6916
rect 41288 6876 41294 6888
rect 33778 6808 33784 6860
rect 33836 6848 33842 6860
rect 34057 6851 34115 6857
rect 33836 6820 33881 6848
rect 33836 6808 33842 6820
rect 34057 6817 34069 6851
rect 34103 6848 34115 6851
rect 34882 6848 34888 6860
rect 34103 6820 34888 6848
rect 34103 6817 34115 6820
rect 34057 6811 34115 6817
rect 34882 6808 34888 6820
rect 34940 6808 34946 6860
rect 35526 6808 35532 6860
rect 35584 6848 35590 6860
rect 35805 6851 35863 6857
rect 35805 6848 35817 6851
rect 35584 6820 35817 6848
rect 35584 6808 35590 6820
rect 35805 6817 35817 6820
rect 35851 6817 35863 6851
rect 35986 6848 35992 6860
rect 35947 6820 35992 6848
rect 35805 6811 35863 6817
rect 35986 6808 35992 6820
rect 36044 6808 36050 6860
rect 36170 6848 36176 6860
rect 36131 6820 36176 6848
rect 36170 6808 36176 6820
rect 36228 6808 36234 6860
rect 36354 6848 36360 6860
rect 36315 6820 36360 6848
rect 36354 6808 36360 6820
rect 36412 6808 36418 6860
rect 36446 6808 36452 6860
rect 36504 6848 36510 6860
rect 36633 6851 36691 6857
rect 36633 6848 36645 6851
rect 36504 6820 36645 6848
rect 36504 6808 36510 6820
rect 36633 6817 36645 6820
rect 36679 6848 36691 6851
rect 36998 6848 37004 6860
rect 36679 6820 37004 6848
rect 36679 6817 36691 6820
rect 36633 6811 36691 6817
rect 36998 6808 37004 6820
rect 37056 6848 37062 6860
rect 37550 6848 37556 6860
rect 37056 6820 37556 6848
rect 37056 6808 37062 6820
rect 37550 6808 37556 6820
rect 37608 6808 37614 6860
rect 37734 6848 37740 6860
rect 37647 6820 37740 6848
rect 37734 6808 37740 6820
rect 37792 6848 37798 6860
rect 38194 6848 38200 6860
rect 37792 6820 38200 6848
rect 37792 6808 37798 6820
rect 38194 6808 38200 6820
rect 38252 6808 38258 6860
rect 38746 6848 38752 6860
rect 38707 6820 38752 6848
rect 38746 6808 38752 6820
rect 38804 6808 38810 6860
rect 38930 6848 38936 6860
rect 38891 6820 38936 6848
rect 38930 6808 38936 6820
rect 38988 6808 38994 6860
rect 39301 6851 39359 6857
rect 39301 6817 39313 6851
rect 39347 6848 39359 6851
rect 40313 6851 40371 6857
rect 40313 6848 40325 6851
rect 39347 6820 40325 6848
rect 39347 6817 39359 6820
rect 39301 6811 39359 6817
rect 40313 6817 40325 6820
rect 40359 6817 40371 6851
rect 40313 6811 40371 6817
rect 40402 6808 40408 6860
rect 40460 6848 40466 6860
rect 40862 6848 40868 6860
rect 40460 6820 40505 6848
rect 40823 6820 40868 6848
rect 40460 6808 40466 6820
rect 40862 6808 40868 6820
rect 40920 6808 40926 6860
rect 41877 6851 41935 6857
rect 41877 6817 41889 6851
rect 41923 6817 41935 6851
rect 41877 6811 41935 6817
rect 29840 6752 32720 6780
rect 33152 6752 33732 6780
rect 35345 6783 35403 6789
rect 27580 6684 28120 6712
rect 31113 6715 31171 6721
rect 27580 6672 27586 6684
rect 31113 6681 31125 6715
rect 31159 6712 31171 6715
rect 32490 6712 32496 6724
rect 31159 6684 32496 6712
rect 31159 6681 31171 6684
rect 31113 6675 31171 6681
rect 32490 6672 32496 6684
rect 32548 6672 32554 6724
rect 32858 6712 32864 6724
rect 32819 6684 32864 6712
rect 32858 6672 32864 6684
rect 32916 6672 32922 6724
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 5592 6616 6837 6644
rect 5592 6604 5598 6616
rect 6825 6613 6837 6616
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 10226 6604 10232 6656
rect 10284 6644 10290 6656
rect 13078 6644 13084 6656
rect 10284 6616 13084 6644
rect 10284 6604 10290 6616
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 14090 6644 14096 6656
rect 14051 6616 14096 6644
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 20254 6644 20260 6656
rect 19392 6616 20260 6644
rect 19392 6604 19398 6616
rect 20254 6604 20260 6616
rect 20312 6604 20318 6656
rect 26602 6604 26608 6656
rect 26660 6644 26666 6656
rect 29454 6644 29460 6656
rect 26660 6616 29460 6644
rect 26660 6604 26666 6616
rect 29454 6604 29460 6616
rect 29512 6604 29518 6656
rect 30006 6644 30012 6656
rect 29967 6616 30012 6644
rect 30006 6604 30012 6616
rect 30064 6604 30070 6656
rect 30098 6604 30104 6656
rect 30156 6644 30162 6656
rect 33152 6644 33180 6752
rect 35345 6749 35357 6783
rect 35391 6780 35403 6783
rect 40129 6783 40187 6789
rect 40129 6780 40141 6783
rect 35391 6752 40141 6780
rect 35391 6749 35403 6752
rect 35345 6743 35403 6749
rect 40129 6749 40141 6752
rect 40175 6780 40187 6783
rect 41598 6780 41604 6792
rect 40175 6752 41604 6780
rect 40175 6749 40187 6752
rect 40129 6743 40187 6749
rect 41598 6740 41604 6752
rect 41656 6780 41662 6792
rect 41693 6783 41751 6789
rect 41693 6780 41705 6783
rect 41656 6752 41705 6780
rect 41656 6740 41662 6752
rect 41693 6749 41705 6752
rect 41739 6749 41751 6783
rect 41892 6780 41920 6811
rect 41966 6808 41972 6860
rect 42024 6848 42030 6860
rect 42024 6820 42069 6848
rect 42168 6820 42656 6848
rect 42024 6808 42030 6820
rect 42168 6780 42196 6820
rect 41892 6752 42196 6780
rect 42429 6783 42487 6789
rect 41693 6743 41751 6749
rect 42429 6749 42441 6783
rect 42475 6749 42487 6783
rect 42628 6780 42656 6820
rect 42702 6808 42708 6860
rect 42760 6848 42766 6860
rect 43349 6851 43407 6857
rect 43349 6848 43361 6851
rect 42760 6820 43361 6848
rect 42760 6808 42766 6820
rect 43349 6817 43361 6820
rect 43395 6817 43407 6851
rect 43898 6848 43904 6860
rect 43859 6820 43904 6848
rect 43349 6811 43407 6817
rect 43898 6808 43904 6820
rect 43956 6808 43962 6860
rect 44177 6851 44235 6857
rect 44177 6817 44189 6851
rect 44223 6848 44235 6851
rect 44266 6848 44272 6860
rect 44223 6820 44272 6848
rect 44223 6817 44235 6820
rect 44177 6811 44235 6817
rect 44266 6808 44272 6820
rect 44324 6808 44330 6860
rect 45189 6851 45247 6857
rect 45189 6817 45201 6851
rect 45235 6817 45247 6851
rect 45189 6811 45247 6817
rect 45465 6851 45523 6857
rect 45465 6817 45477 6851
rect 45511 6848 45523 6851
rect 45646 6848 45652 6860
rect 45511 6820 45652 6848
rect 45511 6817 45523 6820
rect 45465 6811 45523 6817
rect 43438 6780 43444 6792
rect 42628 6752 43444 6780
rect 42429 6743 42487 6749
rect 33318 6672 33324 6724
rect 33376 6712 33382 6724
rect 33873 6715 33931 6721
rect 33873 6712 33885 6715
rect 33376 6684 33885 6712
rect 33376 6672 33382 6684
rect 33873 6681 33885 6684
rect 33919 6712 33931 6715
rect 41046 6712 41052 6724
rect 33919 6684 41052 6712
rect 33919 6681 33931 6684
rect 33873 6675 33931 6681
rect 41046 6672 41052 6684
rect 41104 6672 41110 6724
rect 42444 6712 42472 6743
rect 43438 6740 43444 6752
rect 43496 6740 43502 6792
rect 44358 6780 44364 6792
rect 44319 6752 44364 6780
rect 44358 6740 44364 6752
rect 44416 6780 44422 6792
rect 44910 6780 44916 6792
rect 44416 6752 44916 6780
rect 44416 6740 44422 6752
rect 44910 6740 44916 6752
rect 44968 6740 44974 6792
rect 45204 6780 45232 6811
rect 45646 6808 45652 6820
rect 45704 6808 45710 6860
rect 46750 6848 46756 6860
rect 46711 6820 46756 6848
rect 46750 6808 46756 6820
rect 46808 6808 46814 6860
rect 47026 6848 47032 6860
rect 46987 6820 47032 6848
rect 47026 6808 47032 6820
rect 47084 6808 47090 6860
rect 51092 6857 51120 6888
rect 51350 6876 51356 6888
rect 51408 6876 51414 6928
rect 52457 6919 52515 6925
rect 52457 6885 52469 6919
rect 52503 6916 52515 6919
rect 52546 6916 52552 6928
rect 52503 6888 52552 6916
rect 52503 6885 52515 6888
rect 52457 6879 52515 6885
rect 52546 6876 52552 6888
rect 52604 6876 52610 6928
rect 53190 6916 53196 6928
rect 53116 6888 53196 6916
rect 49053 6851 49111 6857
rect 49053 6848 49065 6851
rect 47136 6820 49065 6848
rect 46106 6780 46112 6792
rect 45204 6752 46112 6780
rect 46106 6740 46112 6752
rect 46164 6740 46170 6792
rect 46566 6740 46572 6792
rect 46624 6780 46630 6792
rect 47136 6780 47164 6820
rect 49053 6817 49065 6820
rect 49099 6817 49111 6851
rect 49053 6811 49111 6817
rect 51077 6851 51135 6857
rect 51077 6817 51089 6851
rect 51123 6817 51135 6851
rect 51077 6811 51135 6817
rect 51169 6851 51227 6857
rect 51169 6817 51181 6851
rect 51215 6848 51227 6851
rect 51258 6848 51264 6860
rect 51215 6820 51264 6848
rect 51215 6817 51227 6820
rect 51169 6811 51227 6817
rect 47302 6780 47308 6792
rect 46624 6752 47164 6780
rect 47263 6752 47308 6780
rect 46624 6740 46630 6752
rect 47302 6740 47308 6752
rect 47360 6740 47366 6792
rect 48682 6740 48688 6792
rect 48740 6780 48746 6792
rect 48961 6783 49019 6789
rect 48961 6780 48973 6783
rect 48740 6752 48973 6780
rect 48740 6740 48746 6752
rect 48961 6749 48973 6752
rect 49007 6749 49019 6783
rect 49068 6780 49096 6811
rect 51258 6808 51264 6820
rect 51316 6808 51322 6860
rect 53116 6857 53144 6888
rect 53190 6876 53196 6888
rect 53248 6876 53254 6928
rect 53650 6876 53656 6928
rect 53708 6916 53714 6928
rect 53708 6888 55076 6916
rect 53708 6876 53714 6888
rect 53101 6851 53159 6857
rect 53101 6817 53113 6851
rect 53147 6817 53159 6851
rect 53101 6811 53159 6817
rect 53469 6851 53527 6857
rect 53469 6817 53481 6851
rect 53515 6848 53527 6851
rect 53834 6848 53840 6860
rect 53515 6820 53840 6848
rect 53515 6817 53527 6820
rect 53469 6811 53527 6817
rect 49326 6780 49332 6792
rect 49068 6752 49332 6780
rect 48961 6743 49019 6749
rect 49326 6740 49332 6752
rect 49384 6740 49390 6792
rect 49510 6780 49516 6792
rect 49471 6752 49516 6780
rect 49510 6740 49516 6752
rect 49568 6740 49574 6792
rect 52362 6780 52368 6792
rect 51000 6752 52368 6780
rect 45281 6715 45339 6721
rect 45281 6712 45293 6715
rect 42444 6684 45293 6712
rect 45281 6681 45293 6684
rect 45327 6681 45339 6715
rect 46842 6712 46848 6724
rect 46803 6684 46848 6712
rect 45281 6675 45339 6681
rect 46842 6672 46848 6684
rect 46900 6672 46906 6724
rect 51000 6712 51028 6752
rect 52362 6740 52368 6752
rect 52420 6740 52426 6792
rect 53193 6783 53251 6789
rect 53193 6749 53205 6783
rect 53239 6780 53251 6783
rect 53282 6780 53288 6792
rect 53239 6752 53288 6780
rect 53239 6749 53251 6752
rect 53193 6743 53251 6749
rect 53282 6740 53288 6752
rect 53340 6740 53346 6792
rect 46952 6684 51028 6712
rect 30156 6616 33180 6644
rect 30156 6604 30162 6616
rect 33226 6604 33232 6656
rect 33284 6644 33290 6656
rect 39482 6644 39488 6656
rect 33284 6616 39488 6644
rect 33284 6604 33290 6616
rect 39482 6604 39488 6616
rect 39540 6604 39546 6656
rect 42610 6604 42616 6656
rect 42668 6644 42674 6656
rect 46952 6644 46980 6684
rect 52178 6672 52184 6724
rect 52236 6712 52242 6724
rect 53484 6712 53512 6811
rect 53834 6808 53840 6820
rect 53892 6808 53898 6860
rect 54754 6848 54760 6860
rect 54715 6820 54760 6848
rect 54754 6808 54760 6820
rect 54812 6808 54818 6860
rect 54941 6851 54999 6857
rect 54941 6817 54953 6851
rect 54987 6817 54999 6851
rect 55048 6848 55076 6888
rect 56134 6848 56140 6860
rect 55048 6820 56140 6848
rect 54941 6811 54999 6817
rect 53561 6783 53619 6789
rect 53561 6749 53573 6783
rect 53607 6749 53619 6783
rect 53561 6743 53619 6749
rect 52236 6684 53512 6712
rect 52236 6672 52242 6684
rect 42668 6616 46980 6644
rect 42668 6604 42674 6616
rect 47026 6604 47032 6656
rect 47084 6644 47090 6656
rect 47946 6644 47952 6656
rect 47084 6616 47952 6644
rect 47084 6604 47090 6616
rect 47946 6604 47952 6616
rect 48004 6604 48010 6656
rect 48038 6604 48044 6656
rect 48096 6644 48102 6656
rect 51258 6644 51264 6656
rect 48096 6616 51264 6644
rect 48096 6604 48102 6616
rect 51258 6604 51264 6616
rect 51316 6604 51322 6656
rect 51353 6647 51411 6653
rect 51353 6613 51365 6647
rect 51399 6644 51411 6647
rect 52914 6644 52920 6656
rect 51399 6616 52920 6644
rect 51399 6613 51411 6616
rect 51353 6607 51411 6613
rect 52914 6604 52920 6616
rect 52972 6604 52978 6656
rect 53006 6604 53012 6656
rect 53064 6644 53070 6656
rect 53576 6644 53604 6743
rect 53742 6740 53748 6792
rect 53800 6780 53806 6792
rect 54956 6780 54984 6811
rect 56134 6808 56140 6820
rect 56192 6808 56198 6860
rect 56686 6848 56692 6860
rect 56647 6820 56692 6848
rect 56686 6808 56692 6820
rect 56744 6808 56750 6860
rect 56796 6848 56824 6956
rect 58069 6919 58127 6925
rect 58069 6885 58081 6919
rect 58115 6916 58127 6919
rect 58618 6916 58624 6928
rect 58115 6888 58624 6916
rect 58115 6885 58127 6888
rect 58069 6879 58127 6885
rect 58618 6876 58624 6888
rect 58676 6876 58682 6928
rect 59354 6876 59360 6928
rect 59412 6916 59418 6928
rect 60737 6919 60795 6925
rect 60737 6916 60749 6919
rect 59412 6888 60749 6916
rect 59412 6876 59418 6888
rect 60737 6885 60749 6888
rect 60783 6885 60795 6919
rect 60737 6879 60795 6885
rect 56962 6848 56968 6860
rect 56796 6820 56968 6848
rect 56962 6808 56968 6820
rect 57020 6808 57026 6860
rect 57241 6851 57299 6857
rect 57241 6817 57253 6851
rect 57287 6848 57299 6851
rect 57974 6848 57980 6860
rect 57287 6820 57980 6848
rect 57287 6817 57299 6820
rect 57241 6811 57299 6817
rect 57974 6808 57980 6820
rect 58032 6808 58038 6860
rect 58710 6848 58716 6860
rect 58671 6820 58716 6848
rect 58710 6808 58716 6820
rect 58768 6808 58774 6860
rect 58802 6808 58808 6860
rect 58860 6848 58866 6860
rect 59081 6851 59139 6857
rect 58860 6820 58905 6848
rect 58860 6808 58866 6820
rect 59081 6817 59093 6851
rect 59127 6848 59139 6851
rect 59906 6848 59912 6860
rect 59127 6820 59912 6848
rect 59127 6817 59139 6820
rect 59081 6811 59139 6817
rect 53800 6752 54984 6780
rect 55309 6783 55367 6789
rect 53800 6740 53806 6752
rect 55309 6749 55321 6783
rect 55355 6749 55367 6783
rect 56226 6780 56232 6792
rect 56187 6752 56232 6780
rect 55309 6743 55367 6749
rect 55324 6712 55352 6743
rect 56226 6740 56232 6752
rect 56284 6780 56290 6792
rect 59096 6780 59124 6811
rect 59906 6808 59912 6820
rect 59964 6808 59970 6860
rect 60274 6848 60280 6860
rect 60235 6820 60280 6848
rect 60274 6808 60280 6820
rect 60332 6808 60338 6860
rect 56284 6752 59124 6780
rect 59173 6783 59231 6789
rect 56284 6740 56290 6752
rect 59173 6749 59185 6783
rect 59219 6780 59231 6783
rect 59538 6780 59544 6792
rect 59219 6752 59544 6780
rect 59219 6749 59231 6752
rect 59173 6743 59231 6749
rect 59538 6740 59544 6752
rect 59596 6740 59602 6792
rect 60182 6780 60188 6792
rect 60143 6752 60188 6780
rect 60182 6740 60188 6752
rect 60240 6740 60246 6792
rect 59262 6712 59268 6724
rect 55324 6684 59268 6712
rect 59262 6672 59268 6684
rect 59320 6672 59326 6724
rect 53064 6616 53604 6644
rect 53064 6604 53070 6616
rect 54018 6604 54024 6656
rect 54076 6644 54082 6656
rect 60274 6644 60280 6656
rect 54076 6616 60280 6644
rect 54076 6604 54082 6616
rect 60274 6604 60280 6616
rect 60332 6604 60338 6656
rect 1104 6554 62192 6576
rect 1104 6502 11163 6554
rect 11215 6502 11227 6554
rect 11279 6502 11291 6554
rect 11343 6502 11355 6554
rect 11407 6502 31526 6554
rect 31578 6502 31590 6554
rect 31642 6502 31654 6554
rect 31706 6502 31718 6554
rect 31770 6502 51888 6554
rect 51940 6502 51952 6554
rect 52004 6502 52016 6554
rect 52068 6502 52080 6554
rect 52132 6502 62192 6554
rect 1104 6480 62192 6502
rect 9674 6440 9680 6452
rect 9635 6412 9680 6440
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 23566 6440 23572 6452
rect 13740 6412 23572 6440
rect 13740 6372 13768 6412
rect 23566 6400 23572 6412
rect 23624 6400 23630 6452
rect 28169 6443 28227 6449
rect 28169 6440 28181 6443
rect 27908 6412 28181 6440
rect 6288 6344 13768 6372
rect 16485 6375 16543 6381
rect 3142 6264 3148 6316
rect 3200 6304 3206 6316
rect 3697 6307 3755 6313
rect 3697 6304 3709 6307
rect 3200 6276 3709 6304
rect 3200 6264 3206 6276
rect 3697 6273 3709 6276
rect 3743 6273 3755 6307
rect 5626 6304 5632 6316
rect 3697 6267 3755 6273
rect 4172 6276 5632 6304
rect 2682 6236 2688 6248
rect 2643 6208 2688 6236
rect 2682 6196 2688 6208
rect 2740 6196 2746 6248
rect 4172 6245 4200 6276
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6205 4215 6239
rect 4157 6199 4215 6205
rect 4430 6196 4436 6248
rect 4488 6236 4494 6248
rect 4525 6239 4583 6245
rect 4525 6236 4537 6239
rect 4488 6208 4537 6236
rect 4488 6196 4494 6208
rect 4525 6205 4537 6208
rect 4571 6205 4583 6239
rect 4525 6199 4583 6205
rect 4617 6239 4675 6245
rect 4617 6205 4629 6239
rect 4663 6236 4675 6239
rect 4798 6236 4804 6248
rect 4663 6208 4804 6236
rect 4663 6205 4675 6208
rect 4617 6199 4675 6205
rect 4798 6196 4804 6208
rect 4856 6236 4862 6248
rect 5350 6236 5356 6248
rect 4856 6208 5356 6236
rect 4856 6196 4862 6208
rect 5350 6196 5356 6208
rect 5408 6236 5414 6248
rect 6288 6236 6316 6344
rect 16485 6341 16497 6375
rect 16531 6372 16543 6375
rect 17126 6372 17132 6384
rect 16531 6344 17132 6372
rect 16531 6341 16543 6344
rect 16485 6335 16543 6341
rect 17126 6332 17132 6344
rect 17184 6332 17190 6384
rect 19886 6372 19892 6384
rect 18064 6344 19892 6372
rect 6362 6264 6368 6316
rect 6420 6304 6426 6316
rect 10134 6304 10140 6316
rect 6420 6276 8248 6304
rect 10095 6276 10140 6304
rect 6420 6264 6426 6276
rect 5408 6208 6316 6236
rect 5408 6196 5414 6208
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 8220 6245 8248 6276
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 10689 6307 10747 6313
rect 10689 6273 10701 6307
rect 10735 6304 10747 6307
rect 11974 6304 11980 6316
rect 10735 6276 11980 6304
rect 10735 6273 10747 6276
rect 10689 6267 10747 6273
rect 11974 6264 11980 6276
rect 12032 6264 12038 6316
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 12526 6304 12532 6316
rect 12483 6276 12532 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 12526 6264 12532 6276
rect 12584 6304 12590 6316
rect 16206 6304 16212 6316
rect 12584 6276 16212 6304
rect 12584 6264 12590 6276
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 16298 6264 16304 6316
rect 16356 6304 16362 6316
rect 16945 6307 17003 6313
rect 16945 6304 16957 6307
rect 16356 6276 16957 6304
rect 16356 6264 16362 6276
rect 16945 6273 16957 6276
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6972 6208 7021 6236
rect 6972 6196 6978 6208
rect 7009 6205 7021 6208
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6205 8263 6239
rect 10226 6236 10232 6248
rect 10187 6208 10232 6236
rect 8205 6199 8263 6205
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 10594 6236 10600 6248
rect 10555 6208 10600 6236
rect 10594 6196 10600 6208
rect 10652 6196 10658 6248
rect 13173 6239 13231 6245
rect 13173 6205 13185 6239
rect 13219 6236 13231 6239
rect 15197 6239 15255 6245
rect 13219 6208 15148 6236
rect 13219 6205 13231 6208
rect 13173 6199 13231 6205
rect 6825 6171 6883 6177
rect 6825 6137 6837 6171
rect 6871 6137 6883 6171
rect 6825 6131 6883 6137
rect 2774 6060 2780 6112
rect 2832 6100 2838 6112
rect 6840 6100 6868 6131
rect 12526 6128 12532 6180
rect 12584 6168 12590 6180
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 12584 6140 12817 6168
rect 12584 6128 12590 6140
rect 12805 6137 12817 6140
rect 12851 6137 12863 6171
rect 15010 6168 15016 6180
rect 14971 6140 15016 6168
rect 12805 6131 12863 6137
rect 15010 6128 15016 6140
rect 15068 6128 15074 6180
rect 15120 6168 15148 6208
rect 15197 6205 15209 6239
rect 15243 6236 15255 6239
rect 15470 6236 15476 6248
rect 15243 6208 15476 6236
rect 15243 6205 15255 6208
rect 15197 6199 15255 6205
rect 15470 6196 15476 6208
rect 15528 6196 15534 6248
rect 16393 6239 16451 6245
rect 16393 6205 16405 6239
rect 16439 6236 16451 6239
rect 16574 6236 16580 6248
rect 16439 6208 16580 6236
rect 16439 6205 16451 6208
rect 16393 6199 16451 6205
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 18064 6245 18092 6344
rect 19886 6332 19892 6344
rect 19944 6372 19950 6384
rect 20070 6372 20076 6384
rect 19944 6344 20076 6372
rect 19944 6332 19950 6344
rect 20070 6332 20076 6344
rect 20128 6332 20134 6384
rect 20162 6332 20168 6384
rect 20220 6372 20226 6384
rect 21361 6375 21419 6381
rect 21361 6372 21373 6375
rect 20220 6344 21373 6372
rect 20220 6332 20226 6344
rect 21361 6341 21373 6344
rect 21407 6341 21419 6375
rect 21361 6335 21419 6341
rect 19518 6304 19524 6316
rect 19479 6276 19524 6304
rect 19518 6264 19524 6276
rect 19576 6264 19582 6316
rect 20714 6304 20720 6316
rect 20088 6276 20720 6304
rect 16669 6239 16727 6245
rect 16669 6205 16681 6239
rect 16715 6236 16727 6239
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 16715 6208 18061 6236
rect 16715 6205 16727 6208
rect 16669 6199 16727 6205
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 19429 6239 19487 6245
rect 19429 6205 19441 6239
rect 19475 6236 19487 6239
rect 20088 6236 20116 6276
rect 20714 6264 20720 6276
rect 20772 6264 20778 6316
rect 21376 6304 21404 6335
rect 27798 6332 27804 6384
rect 27856 6372 27862 6384
rect 27908 6372 27936 6412
rect 28169 6409 28181 6412
rect 28215 6409 28227 6443
rect 28169 6403 28227 6409
rect 28258 6400 28264 6452
rect 28316 6440 28322 6452
rect 33226 6440 33232 6452
rect 28316 6412 33232 6440
rect 28316 6400 28322 6412
rect 33226 6400 33232 6412
rect 33284 6400 33290 6452
rect 36170 6440 36176 6452
rect 33336 6412 36176 6440
rect 27856 6344 27936 6372
rect 27856 6332 27862 6344
rect 28350 6332 28356 6384
rect 28408 6372 28414 6384
rect 33336 6372 33364 6412
rect 36170 6400 36176 6412
rect 36228 6440 36234 6452
rect 36906 6440 36912 6452
rect 36228 6412 36912 6440
rect 36228 6400 36234 6412
rect 36906 6400 36912 6412
rect 36964 6400 36970 6452
rect 38838 6400 38844 6452
rect 38896 6440 38902 6452
rect 40678 6440 40684 6452
rect 38896 6412 40684 6440
rect 38896 6400 38902 6412
rect 40678 6400 40684 6412
rect 40736 6400 40742 6452
rect 40773 6443 40831 6449
rect 40773 6409 40785 6443
rect 40819 6440 40831 6443
rect 41966 6440 41972 6452
rect 40819 6412 41972 6440
rect 40819 6409 40831 6412
rect 40773 6403 40831 6409
rect 41966 6400 41972 6412
rect 42024 6400 42030 6452
rect 42334 6400 42340 6452
rect 42392 6440 42398 6452
rect 48314 6440 48320 6452
rect 42392 6412 48320 6440
rect 42392 6400 42398 6412
rect 48314 6400 48320 6412
rect 48372 6400 48378 6452
rect 53006 6440 53012 6452
rect 49712 6412 53012 6440
rect 28408 6344 33364 6372
rect 28408 6332 28414 6344
rect 35986 6332 35992 6384
rect 36044 6372 36050 6384
rect 36446 6372 36452 6384
rect 36044 6344 36452 6372
rect 36044 6332 36050 6344
rect 36446 6332 36452 6344
rect 36504 6332 36510 6384
rect 36814 6332 36820 6384
rect 36872 6372 36878 6384
rect 38930 6372 38936 6384
rect 36872 6344 38936 6372
rect 36872 6332 36878 6344
rect 38930 6332 38936 6344
rect 38988 6332 38994 6384
rect 39666 6332 39672 6384
rect 39724 6372 39730 6384
rect 49326 6372 49332 6384
rect 39724 6344 49332 6372
rect 39724 6332 39730 6344
rect 49326 6332 49332 6344
rect 49384 6332 49390 6384
rect 25222 6304 25228 6316
rect 21376 6276 25084 6304
rect 25183 6276 25228 6304
rect 20254 6236 20260 6248
rect 19475 6208 20116 6236
rect 20215 6208 20260 6236
rect 19475 6205 19487 6208
rect 19429 6199 19487 6205
rect 20254 6196 20260 6208
rect 20312 6196 20318 6248
rect 20346 6196 20352 6248
rect 20404 6236 20410 6248
rect 20404 6208 20449 6236
rect 20404 6196 20410 6208
rect 20806 6196 20812 6248
rect 20864 6236 20870 6248
rect 21269 6239 21327 6245
rect 21269 6236 21281 6239
rect 20864 6208 21281 6236
rect 20864 6196 20870 6208
rect 21269 6205 21281 6208
rect 21315 6205 21327 6239
rect 21542 6236 21548 6248
rect 21503 6208 21548 6236
rect 21269 6199 21327 6205
rect 21542 6196 21548 6208
rect 21600 6196 21606 6248
rect 21910 6196 21916 6248
rect 21968 6236 21974 6248
rect 23845 6239 23903 6245
rect 23845 6236 23857 6239
rect 21968 6208 23857 6236
rect 21968 6196 21974 6208
rect 23845 6205 23857 6208
rect 23891 6236 23903 6239
rect 24946 6236 24952 6248
rect 23891 6208 24164 6236
rect 24907 6208 24952 6236
rect 23891 6205 23903 6208
rect 23845 6199 23903 6205
rect 22738 6168 22744 6180
rect 15120 6140 22744 6168
rect 22738 6128 22744 6140
rect 22796 6128 22802 6180
rect 7006 6100 7012 6112
rect 2832 6072 2877 6100
rect 6840 6072 7012 6100
rect 2832 6060 2838 6072
rect 7006 6060 7012 6072
rect 7064 6060 7070 6112
rect 7098 6060 7104 6112
rect 7156 6100 7162 6112
rect 7156 6072 7201 6100
rect 7156 6060 7162 6072
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 8297 6103 8355 6109
rect 8297 6100 8309 6103
rect 7340 6072 8309 6100
rect 7340 6060 7346 6072
rect 8297 6069 8309 6072
rect 8343 6069 8355 6103
rect 8297 6063 8355 6069
rect 12066 6060 12072 6112
rect 12124 6100 12130 6112
rect 12618 6100 12624 6112
rect 12124 6072 12624 6100
rect 12124 6060 12130 6072
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 15289 6103 15347 6109
rect 12768 6072 12813 6100
rect 12768 6060 12774 6072
rect 15289 6069 15301 6103
rect 15335 6100 15347 6103
rect 16666 6100 16672 6112
rect 15335 6072 16672 6100
rect 15335 6069 15347 6072
rect 15289 6063 15347 6069
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 18233 6103 18291 6109
rect 18233 6069 18245 6103
rect 18279 6100 18291 6103
rect 18690 6100 18696 6112
rect 18279 6072 18696 6100
rect 18279 6069 18291 6072
rect 18233 6063 18291 6069
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 21726 6100 21732 6112
rect 21687 6072 21732 6100
rect 21726 6060 21732 6072
rect 21784 6060 21790 6112
rect 24026 6100 24032 6112
rect 23987 6072 24032 6100
rect 24026 6060 24032 6072
rect 24084 6060 24090 6112
rect 24136 6100 24164 6208
rect 24946 6196 24952 6208
rect 25004 6196 25010 6248
rect 25056 6236 25084 6276
rect 25222 6264 25228 6276
rect 25280 6264 25286 6316
rect 31435 6307 31493 6313
rect 31435 6304 31447 6307
rect 27908 6276 31447 6304
rect 27908 6236 27936 6276
rect 31435 6273 31447 6276
rect 31481 6304 31493 6307
rect 33318 6304 33324 6316
rect 31481 6276 33324 6304
rect 31481 6273 31493 6276
rect 31435 6267 31493 6273
rect 33318 6264 33324 6276
rect 33376 6264 33382 6316
rect 39025 6307 39083 6313
rect 39025 6304 39037 6307
rect 33520 6276 39037 6304
rect 25056 6208 27936 6236
rect 27985 6239 28043 6245
rect 27985 6205 27997 6239
rect 28031 6236 28043 6239
rect 28902 6236 28908 6248
rect 28031 6208 28908 6236
rect 28031 6205 28043 6208
rect 27985 6199 28043 6205
rect 28902 6196 28908 6208
rect 28960 6196 28966 6248
rect 29273 6239 29331 6245
rect 29273 6205 29285 6239
rect 29319 6236 29331 6239
rect 29362 6236 29368 6248
rect 29319 6208 29368 6236
rect 29319 6205 29331 6208
rect 29273 6199 29331 6205
rect 29362 6196 29368 6208
rect 29420 6196 29426 6248
rect 29454 6196 29460 6248
rect 29512 6236 29518 6248
rect 31202 6236 31208 6248
rect 29512 6208 31208 6236
rect 29512 6196 29518 6208
rect 31202 6196 31208 6208
rect 31260 6196 31266 6248
rect 31294 6196 31300 6248
rect 31352 6236 31358 6248
rect 31573 6239 31631 6245
rect 31352 6208 31397 6236
rect 31352 6196 31358 6208
rect 31573 6205 31585 6239
rect 31619 6205 31631 6239
rect 31573 6199 31631 6205
rect 25884 6140 30052 6168
rect 25884 6100 25912 6140
rect 30024 6112 30052 6140
rect 30466 6128 30472 6180
rect 30524 6168 30530 6180
rect 30745 6171 30803 6177
rect 30745 6168 30757 6171
rect 30524 6140 30757 6168
rect 30524 6128 30530 6140
rect 30745 6137 30757 6140
rect 30791 6137 30803 6171
rect 30745 6131 30803 6137
rect 30926 6128 30932 6180
rect 30984 6168 30990 6180
rect 31588 6168 31616 6199
rect 31754 6196 31760 6248
rect 31812 6236 31818 6248
rect 33520 6236 33548 6276
rect 39025 6273 39037 6276
rect 39071 6304 39083 6307
rect 39390 6304 39396 6316
rect 39071 6276 39396 6304
rect 39071 6273 39083 6276
rect 39025 6267 39083 6273
rect 39390 6264 39396 6276
rect 39448 6264 39454 6316
rect 39577 6307 39635 6313
rect 39577 6273 39589 6307
rect 39623 6304 39635 6307
rect 41690 6304 41696 6316
rect 39623 6276 41696 6304
rect 39623 6273 39635 6276
rect 39577 6267 39635 6273
rect 41690 6264 41696 6276
rect 41748 6264 41754 6316
rect 44910 6264 44916 6316
rect 44968 6304 44974 6316
rect 47949 6307 48007 6313
rect 44968 6276 46612 6304
rect 44968 6264 44974 6276
rect 31812 6208 33548 6236
rect 33577 6239 33635 6245
rect 31812 6196 31818 6208
rect 33577 6205 33589 6239
rect 33623 6236 33635 6239
rect 34054 6236 34060 6248
rect 33623 6208 34060 6236
rect 33623 6205 33635 6208
rect 33577 6199 33635 6205
rect 34054 6196 34060 6208
rect 34112 6196 34118 6248
rect 34238 6196 34244 6248
rect 34296 6236 34302 6248
rect 34885 6239 34943 6245
rect 34885 6236 34897 6239
rect 34296 6208 34897 6236
rect 34296 6196 34302 6208
rect 34885 6205 34897 6208
rect 34931 6205 34943 6239
rect 34885 6199 34943 6205
rect 36173 6239 36231 6245
rect 36173 6205 36185 6239
rect 36219 6205 36231 6239
rect 36446 6236 36452 6248
rect 36407 6208 36452 6236
rect 36173 6199 36231 6205
rect 30984 6140 31616 6168
rect 33413 6171 33471 6177
rect 30984 6128 30990 6140
rect 33413 6137 33425 6171
rect 33459 6137 33471 6171
rect 33413 6131 33471 6137
rect 33965 6171 34023 6177
rect 33965 6137 33977 6171
rect 34011 6168 34023 6171
rect 35894 6168 35900 6180
rect 34011 6140 35900 6168
rect 34011 6137 34023 6140
rect 33965 6131 34023 6137
rect 24136 6072 25912 6100
rect 25958 6060 25964 6112
rect 26016 6100 26022 6112
rect 26513 6103 26571 6109
rect 26513 6100 26525 6103
rect 26016 6072 26525 6100
rect 26016 6060 26022 6072
rect 26513 6069 26525 6072
rect 26559 6100 26571 6103
rect 29270 6100 29276 6112
rect 26559 6072 29276 6100
rect 26559 6069 26571 6072
rect 26513 6063 26571 6069
rect 29270 6060 29276 6072
rect 29328 6060 29334 6112
rect 29454 6100 29460 6112
rect 29415 6072 29460 6100
rect 29454 6060 29460 6072
rect 29512 6060 29518 6112
rect 30006 6060 30012 6112
rect 30064 6100 30070 6112
rect 33428 6100 33456 6131
rect 35894 6128 35900 6140
rect 35952 6128 35958 6180
rect 35066 6100 35072 6112
rect 30064 6072 33456 6100
rect 35027 6072 35072 6100
rect 30064 6060 30070 6072
rect 35066 6060 35072 6072
rect 35124 6060 35130 6112
rect 36188 6100 36216 6199
rect 36446 6196 36452 6208
rect 36504 6196 36510 6248
rect 36906 6236 36912 6248
rect 36867 6208 36912 6236
rect 36906 6196 36912 6208
rect 36964 6196 36970 6248
rect 37090 6196 37096 6248
rect 37148 6236 37154 6248
rect 37277 6239 37335 6245
rect 37277 6236 37289 6239
rect 37148 6208 37289 6236
rect 37148 6196 37154 6208
rect 37277 6205 37289 6208
rect 37323 6205 37335 6239
rect 37277 6199 37335 6205
rect 37642 6196 37648 6248
rect 37700 6236 37706 6248
rect 37737 6239 37795 6245
rect 37737 6236 37749 6239
rect 37700 6208 37749 6236
rect 37700 6196 37706 6208
rect 37737 6205 37749 6208
rect 37783 6205 37795 6239
rect 39114 6236 39120 6248
rect 39075 6208 39120 6236
rect 37737 6199 37795 6205
rect 39114 6196 39120 6208
rect 39172 6236 39178 6248
rect 39172 6208 40632 6236
rect 39172 6196 39178 6208
rect 36354 6168 36360 6180
rect 36315 6140 36360 6168
rect 36354 6128 36360 6140
rect 36412 6128 36418 6180
rect 39482 6128 39488 6180
rect 39540 6168 39546 6180
rect 40402 6168 40408 6180
rect 39540 6140 40408 6168
rect 39540 6128 39546 6140
rect 40402 6128 40408 6140
rect 40460 6168 40466 6180
rect 40497 6171 40555 6177
rect 40497 6168 40509 6171
rect 40460 6140 40509 6168
rect 40460 6128 40466 6140
rect 40497 6137 40509 6140
rect 40543 6137 40555 6171
rect 40604 6168 40632 6208
rect 40678 6196 40684 6248
rect 40736 6236 40742 6248
rect 40736 6208 40781 6236
rect 40736 6196 40742 6208
rect 41414 6196 41420 6248
rect 41472 6236 41478 6248
rect 41877 6239 41935 6245
rect 41877 6236 41889 6239
rect 41472 6208 41889 6236
rect 41472 6196 41478 6208
rect 41877 6205 41889 6208
rect 41923 6236 41935 6239
rect 42242 6236 42248 6248
rect 41923 6208 42248 6236
rect 41923 6205 41935 6208
rect 41877 6199 41935 6205
rect 42242 6196 42248 6208
rect 42300 6196 42306 6248
rect 42610 6236 42616 6248
rect 42571 6208 42616 6236
rect 42610 6196 42616 6208
rect 42668 6196 42674 6248
rect 42886 6236 42892 6248
rect 42847 6208 42892 6236
rect 42886 6196 42892 6208
rect 42944 6196 42950 6248
rect 44634 6236 44640 6248
rect 44595 6208 44640 6236
rect 44634 6196 44640 6208
rect 44692 6196 44698 6248
rect 46584 6245 46612 6276
rect 47949 6273 47961 6307
rect 47995 6304 48007 6307
rect 49712 6304 49740 6412
rect 53006 6400 53012 6412
rect 53064 6400 53070 6452
rect 53285 6443 53343 6449
rect 53285 6409 53297 6443
rect 53331 6440 53343 6443
rect 53558 6440 53564 6452
rect 53331 6412 53564 6440
rect 53331 6409 53343 6412
rect 53285 6403 53343 6409
rect 53558 6400 53564 6412
rect 53616 6400 53622 6452
rect 53742 6400 53748 6452
rect 53800 6440 53806 6452
rect 58158 6440 58164 6452
rect 53800 6412 58164 6440
rect 53800 6400 53806 6412
rect 58158 6400 58164 6412
rect 58216 6400 58222 6452
rect 49786 6332 49792 6384
rect 49844 6372 49850 6384
rect 51626 6372 51632 6384
rect 49844 6344 51632 6372
rect 49844 6332 49850 6344
rect 51626 6332 51632 6344
rect 51684 6332 51690 6384
rect 52089 6375 52147 6381
rect 52089 6341 52101 6375
rect 52135 6372 52147 6375
rect 52178 6372 52184 6384
rect 52135 6344 52184 6372
rect 52135 6341 52147 6344
rect 52089 6335 52147 6341
rect 52178 6332 52184 6344
rect 52236 6332 52242 6384
rect 53653 6375 53711 6381
rect 53653 6372 53665 6375
rect 53300 6344 53665 6372
rect 47995 6276 49740 6304
rect 50249 6307 50307 6313
rect 47995 6273 48007 6276
rect 47949 6267 48007 6273
rect 50249 6273 50261 6307
rect 50295 6304 50307 6307
rect 50522 6304 50528 6316
rect 50295 6276 50528 6304
rect 50295 6273 50307 6276
rect 50249 6267 50307 6273
rect 50522 6264 50528 6276
rect 50580 6264 50586 6316
rect 51166 6264 51172 6316
rect 51224 6304 51230 6316
rect 53300 6304 53328 6344
rect 53653 6341 53665 6344
rect 53699 6372 53711 6375
rect 56686 6372 56692 6384
rect 53699 6344 56692 6372
rect 53699 6341 53711 6344
rect 53653 6335 53711 6341
rect 56686 6332 56692 6344
rect 56744 6372 56750 6384
rect 56744 6344 60964 6372
rect 56744 6332 56750 6344
rect 51224 6276 53328 6304
rect 53377 6307 53435 6313
rect 51224 6264 51230 6276
rect 53377 6273 53389 6307
rect 53423 6304 53435 6307
rect 53558 6304 53564 6316
rect 53423 6276 53564 6304
rect 53423 6273 53435 6276
rect 53377 6267 53435 6273
rect 53558 6264 53564 6276
rect 53616 6304 53622 6316
rect 53926 6304 53932 6316
rect 53616 6276 53932 6304
rect 53616 6264 53622 6276
rect 53926 6264 53932 6276
rect 53984 6264 53990 6316
rect 54662 6264 54668 6316
rect 54720 6304 54726 6316
rect 54720 6276 59124 6304
rect 54720 6264 54726 6276
rect 44729 6239 44787 6245
rect 44729 6205 44741 6239
rect 44775 6205 44787 6239
rect 44729 6199 44787 6205
rect 45189 6239 45247 6245
rect 45189 6205 45201 6239
rect 45235 6236 45247 6239
rect 46569 6239 46627 6245
rect 45235 6208 46520 6236
rect 45235 6205 45247 6208
rect 45189 6199 45247 6205
rect 42334 6168 42340 6180
rect 40604 6140 42340 6168
rect 40497 6131 40555 6137
rect 42334 6128 42340 6140
rect 42392 6128 42398 6180
rect 42426 6128 42432 6180
rect 42484 6168 42490 6180
rect 44744 6168 44772 6199
rect 46290 6168 46296 6180
rect 42484 6140 46296 6168
rect 42484 6128 42490 6140
rect 46290 6128 46296 6140
rect 46348 6128 46354 6180
rect 46385 6171 46443 6177
rect 46385 6137 46397 6171
rect 46431 6137 46443 6171
rect 46492 6168 46520 6208
rect 46569 6205 46581 6239
rect 46615 6205 46627 6239
rect 46569 6199 46627 6205
rect 46937 6239 46995 6245
rect 46937 6205 46949 6239
rect 46983 6236 46995 6239
rect 47857 6239 47915 6245
rect 47857 6236 47869 6239
rect 46983 6208 47869 6236
rect 46983 6205 46995 6208
rect 46937 6199 46995 6205
rect 47857 6205 47869 6208
rect 47903 6205 47915 6239
rect 48682 6236 48688 6248
rect 48643 6208 48688 6236
rect 47857 6199 47915 6205
rect 48682 6196 48688 6208
rect 48740 6196 48746 6248
rect 48777 6239 48835 6245
rect 48777 6205 48789 6239
rect 48823 6236 48835 6239
rect 48866 6236 48872 6248
rect 48823 6208 48872 6236
rect 48823 6205 48835 6208
rect 48777 6199 48835 6205
rect 48866 6196 48872 6208
rect 48924 6236 48930 6248
rect 49510 6236 49516 6248
rect 48924 6208 49516 6236
rect 48924 6196 48930 6208
rect 49510 6196 49516 6208
rect 49568 6196 49574 6248
rect 50382 6239 50440 6245
rect 50382 6205 50394 6239
rect 50428 6236 50440 6239
rect 50614 6236 50620 6248
rect 50428 6208 50620 6236
rect 50428 6205 50440 6208
rect 50382 6199 50440 6205
rect 50614 6196 50620 6208
rect 50672 6196 50678 6248
rect 51442 6196 51448 6248
rect 51500 6236 51506 6248
rect 51905 6239 51963 6245
rect 51905 6236 51917 6239
rect 51500 6208 51917 6236
rect 51500 6196 51506 6208
rect 51905 6205 51917 6208
rect 51951 6205 51963 6239
rect 51905 6199 51963 6205
rect 52822 6196 52828 6248
rect 52880 6236 52886 6248
rect 53156 6239 53214 6245
rect 53156 6236 53168 6239
rect 52880 6208 53168 6236
rect 52880 6196 52886 6208
rect 53156 6205 53168 6208
rect 53202 6205 53214 6239
rect 53156 6199 53214 6205
rect 53282 6196 53288 6248
rect 53340 6236 53346 6248
rect 54478 6236 54484 6248
rect 53340 6208 54484 6236
rect 53340 6196 53346 6208
rect 54478 6196 54484 6208
rect 54536 6196 54542 6248
rect 54570 6196 54576 6248
rect 54628 6236 54634 6248
rect 55122 6236 55128 6248
rect 54628 6208 54673 6236
rect 55083 6208 55128 6236
rect 54628 6196 54634 6208
rect 55122 6196 55128 6208
rect 55180 6196 55186 6248
rect 55398 6236 55404 6248
rect 55359 6208 55404 6236
rect 55398 6196 55404 6208
rect 55456 6196 55462 6248
rect 55585 6239 55643 6245
rect 55585 6236 55597 6239
rect 55508 6208 55597 6236
rect 49602 6168 49608 6180
rect 46492 6140 49608 6168
rect 46385 6131 46443 6137
rect 36446 6100 36452 6112
rect 36188 6072 36452 6100
rect 36446 6060 36452 6072
rect 36504 6100 36510 6112
rect 41969 6103 42027 6109
rect 41969 6100 41981 6103
rect 36504 6072 41981 6100
rect 36504 6060 36510 6072
rect 41969 6069 41981 6072
rect 42015 6069 42027 6103
rect 41969 6063 42027 6069
rect 42794 6060 42800 6112
rect 42852 6100 42858 6112
rect 45554 6100 45560 6112
rect 42852 6072 45560 6100
rect 42852 6060 42858 6072
rect 45554 6060 45560 6072
rect 45612 6060 45618 6112
rect 46400 6100 46428 6131
rect 49602 6128 49608 6140
rect 49660 6128 49666 6180
rect 49786 6128 49792 6180
rect 49844 6168 49850 6180
rect 50801 6171 50859 6177
rect 50801 6168 50813 6171
rect 49844 6140 50813 6168
rect 49844 6128 49850 6140
rect 50801 6137 50813 6140
rect 50847 6137 50859 6171
rect 50801 6131 50859 6137
rect 53006 6128 53012 6180
rect 53064 6168 53070 6180
rect 53064 6140 53109 6168
rect 53064 6128 53070 6140
rect 53742 6128 53748 6180
rect 53800 6168 53806 6180
rect 55508 6168 55536 6208
rect 55585 6205 55597 6208
rect 55631 6236 55643 6239
rect 58710 6236 58716 6248
rect 55631 6208 56364 6236
rect 58671 6208 58716 6236
rect 55631 6205 55643 6208
rect 55585 6199 55643 6205
rect 53800 6140 55536 6168
rect 53800 6128 53806 6140
rect 46750 6100 46756 6112
rect 46400 6072 46756 6100
rect 46750 6060 46756 6072
rect 46808 6100 46814 6112
rect 50706 6100 50712 6112
rect 46808 6072 50712 6100
rect 46808 6060 46814 6072
rect 50706 6060 50712 6072
rect 50764 6060 50770 6112
rect 52178 6060 52184 6112
rect 52236 6100 52242 6112
rect 56226 6100 56232 6112
rect 52236 6072 56232 6100
rect 52236 6060 52242 6072
rect 56226 6060 56232 6072
rect 56284 6060 56290 6112
rect 56336 6100 56364 6208
rect 58710 6196 58716 6208
rect 58768 6196 58774 6248
rect 58802 6196 58808 6248
rect 58860 6236 58866 6248
rect 59096 6245 59124 6276
rect 59262 6264 59268 6316
rect 59320 6304 59326 6316
rect 59320 6276 59400 6304
rect 59320 6264 59326 6276
rect 59081 6239 59139 6245
rect 58860 6208 58905 6236
rect 58860 6196 58866 6208
rect 59081 6205 59093 6239
rect 59127 6205 59139 6239
rect 59081 6199 59139 6205
rect 59170 6196 59176 6248
rect 59228 6236 59234 6248
rect 59372 6236 59400 6276
rect 59538 6264 59544 6316
rect 59596 6304 59602 6316
rect 60093 6307 60151 6313
rect 60093 6304 60105 6307
rect 59596 6276 60105 6304
rect 59596 6264 59602 6276
rect 60093 6273 60105 6276
rect 60139 6273 60151 6307
rect 60093 6267 60151 6273
rect 60200 6276 60780 6304
rect 60200 6236 60228 6276
rect 60752 6245 60780 6276
rect 60936 6245 60964 6344
rect 59228 6208 59273 6236
rect 59372 6208 60228 6236
rect 60553 6239 60611 6245
rect 59228 6196 59234 6208
rect 60553 6205 60565 6239
rect 60599 6205 60611 6239
rect 60553 6199 60611 6205
rect 60737 6239 60795 6245
rect 60737 6205 60749 6239
rect 60783 6205 60795 6239
rect 60737 6199 60795 6205
rect 60921 6239 60979 6245
rect 60921 6205 60933 6239
rect 60967 6205 60979 6239
rect 60921 6199 60979 6205
rect 58066 6168 58072 6180
rect 58027 6140 58072 6168
rect 58066 6128 58072 6140
rect 58124 6128 58130 6180
rect 57790 6100 57796 6112
rect 56336 6072 57796 6100
rect 57790 6060 57796 6072
rect 57848 6100 57854 6112
rect 60568 6100 60596 6199
rect 57848 6072 60596 6100
rect 57848 6060 57854 6072
rect 1104 6010 62192 6032
rect 1104 5958 21344 6010
rect 21396 5958 21408 6010
rect 21460 5958 21472 6010
rect 21524 5958 21536 6010
rect 21588 5958 41707 6010
rect 41759 5958 41771 6010
rect 41823 5958 41835 6010
rect 41887 5958 41899 6010
rect 41951 5958 62192 6010
rect 1104 5936 62192 5958
rect 8202 5896 8208 5908
rect 2608 5868 8208 5896
rect 2608 5769 2636 5868
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 12710 5896 12716 5908
rect 8996 5868 12716 5896
rect 8996 5856 9002 5868
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 13814 5856 13820 5908
rect 13872 5896 13878 5908
rect 23198 5896 23204 5908
rect 13872 5868 23204 5896
rect 13872 5856 13878 5868
rect 23198 5856 23204 5868
rect 23256 5896 23262 5908
rect 27154 5896 27160 5908
rect 23256 5868 27160 5896
rect 23256 5856 23262 5868
rect 27154 5856 27160 5868
rect 27212 5856 27218 5908
rect 27246 5856 27252 5908
rect 27304 5896 27310 5908
rect 30926 5896 30932 5908
rect 27304 5868 30932 5896
rect 27304 5856 27310 5868
rect 30926 5856 30932 5868
rect 30984 5856 30990 5908
rect 31294 5856 31300 5908
rect 31352 5896 31358 5908
rect 35066 5896 35072 5908
rect 31352 5868 35072 5896
rect 31352 5856 31358 5868
rect 35066 5856 35072 5868
rect 35124 5896 35130 5908
rect 37553 5899 37611 5905
rect 37553 5896 37565 5899
rect 35124 5868 37565 5896
rect 35124 5856 35130 5868
rect 37553 5865 37565 5868
rect 37599 5865 37611 5899
rect 37553 5859 37611 5865
rect 37918 5856 37924 5908
rect 37976 5896 37982 5908
rect 38289 5899 38347 5905
rect 38289 5896 38301 5899
rect 37976 5868 38301 5896
rect 37976 5856 37982 5868
rect 38289 5865 38301 5868
rect 38335 5896 38347 5899
rect 39022 5896 39028 5908
rect 38335 5868 39028 5896
rect 38335 5865 38347 5868
rect 38289 5859 38347 5865
rect 39022 5856 39028 5868
rect 39080 5856 39086 5908
rect 42794 5896 42800 5908
rect 41340 5868 42800 5896
rect 4157 5831 4215 5837
rect 4157 5797 4169 5831
rect 4203 5828 4215 5831
rect 4338 5828 4344 5840
rect 4203 5800 4344 5828
rect 4203 5797 4215 5800
rect 4157 5791 4215 5797
rect 4338 5788 4344 5800
rect 4396 5788 4402 5840
rect 5534 5828 5540 5840
rect 4632 5800 5540 5828
rect 2593 5763 2651 5769
rect 2593 5729 2605 5763
rect 2639 5729 2651 5763
rect 2593 5723 2651 5729
rect 2685 5763 2743 5769
rect 2685 5729 2697 5763
rect 2731 5760 2743 5763
rect 4246 5760 4252 5772
rect 2731 5732 4252 5760
rect 2731 5729 2743 5732
rect 2685 5723 2743 5729
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 4632 5769 4660 5800
rect 5534 5788 5540 5800
rect 5592 5788 5598 5840
rect 6730 5828 6736 5840
rect 6196 5800 6736 5828
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5729 4675 5763
rect 4798 5760 4804 5772
rect 4759 5732 4804 5760
rect 4617 5723 4675 5729
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 4985 5763 5043 5769
rect 4985 5729 4997 5763
rect 5031 5760 5043 5763
rect 5718 5760 5724 5772
rect 5031 5732 5724 5760
rect 5031 5729 5043 5732
rect 4985 5723 5043 5729
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 6196 5769 6224 5800
rect 6730 5788 6736 5800
rect 6788 5788 6794 5840
rect 15010 5788 15016 5840
rect 15068 5828 15074 5840
rect 21174 5828 21180 5840
rect 15068 5800 16988 5828
rect 15068 5788 15074 5800
rect 6181 5763 6239 5769
rect 6181 5729 6193 5763
rect 6227 5729 6239 5763
rect 6181 5723 6239 5729
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5729 6607 5763
rect 6549 5723 6607 5729
rect 6825 5763 6883 5769
rect 6825 5729 6837 5763
rect 6871 5760 6883 5763
rect 7282 5760 7288 5772
rect 6871 5732 7288 5760
rect 6871 5729 6883 5732
rect 6825 5723 6883 5729
rect 2866 5556 2872 5568
rect 2827 5528 2872 5556
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 6564 5556 6592 5723
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 7926 5760 7932 5772
rect 7887 5732 7932 5760
rect 7926 5720 7932 5732
rect 7984 5720 7990 5772
rect 8018 5720 8024 5772
rect 8076 5760 8082 5772
rect 8205 5763 8263 5769
rect 8205 5760 8217 5763
rect 8076 5732 8217 5760
rect 8076 5720 8082 5732
rect 8205 5729 8217 5732
rect 8251 5729 8263 5763
rect 8205 5723 8263 5729
rect 11057 5763 11115 5769
rect 11057 5729 11069 5763
rect 11103 5760 11115 5763
rect 11790 5760 11796 5772
rect 11103 5732 11796 5760
rect 11103 5729 11115 5732
rect 11057 5723 11115 5729
rect 11790 5720 11796 5732
rect 11848 5760 11854 5772
rect 12342 5760 12348 5772
rect 11848 5732 12348 5760
rect 11848 5720 11854 5732
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 13541 5763 13599 5769
rect 13541 5760 13553 5763
rect 12492 5732 13553 5760
rect 12492 5720 12498 5732
rect 13541 5729 13553 5732
rect 13587 5729 13599 5763
rect 13541 5723 13599 5729
rect 15194 5720 15200 5772
rect 15252 5760 15258 5772
rect 15473 5763 15531 5769
rect 15473 5760 15485 5763
rect 15252 5732 15485 5760
rect 15252 5720 15258 5732
rect 15473 5729 15485 5732
rect 15519 5729 15531 5763
rect 15654 5760 15660 5772
rect 15615 5732 15660 5760
rect 15473 5723 15531 5729
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 15746 5720 15752 5772
rect 15804 5760 15810 5772
rect 16390 5760 16396 5772
rect 15804 5732 16396 5760
rect 15804 5720 15810 5732
rect 16390 5720 16396 5732
rect 16448 5760 16454 5772
rect 16853 5763 16911 5769
rect 16853 5760 16865 5763
rect 16448 5732 16865 5760
rect 16448 5720 16454 5732
rect 16853 5729 16865 5732
rect 16899 5729 16911 5763
rect 16960 5760 16988 5800
rect 19260 5800 21180 5828
rect 19260 5760 19288 5800
rect 21174 5788 21180 5800
rect 21232 5788 21238 5840
rect 23293 5831 23351 5837
rect 23293 5797 23305 5831
rect 23339 5828 23351 5831
rect 23474 5828 23480 5840
rect 23339 5800 23480 5828
rect 23339 5797 23351 5800
rect 23293 5791 23351 5797
rect 23474 5788 23480 5800
rect 23532 5788 23538 5840
rect 25590 5788 25596 5840
rect 25648 5828 25654 5840
rect 26513 5831 26571 5837
rect 26513 5828 26525 5831
rect 25648 5800 26525 5828
rect 25648 5788 25654 5800
rect 26513 5797 26525 5800
rect 26559 5797 26571 5831
rect 27982 5828 27988 5840
rect 26513 5791 26571 5797
rect 26804 5800 27384 5828
rect 16960 5732 19288 5760
rect 16853 5723 16911 5729
rect 19334 5720 19340 5772
rect 19392 5760 19398 5772
rect 19521 5763 19579 5769
rect 19392 5732 19437 5760
rect 19392 5720 19398 5732
rect 19521 5729 19533 5763
rect 19567 5760 19579 5763
rect 21082 5760 21088 5772
rect 19567 5732 21088 5760
rect 19567 5729 19579 5732
rect 19521 5723 19579 5729
rect 21082 5720 21088 5732
rect 21140 5720 21146 5772
rect 23385 5763 23443 5769
rect 23385 5729 23397 5763
rect 23431 5729 23443 5763
rect 24854 5760 24860 5772
rect 24815 5732 24860 5760
rect 23385 5723 23443 5729
rect 8386 5692 8392 5704
rect 8347 5664 8392 5692
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 11333 5695 11391 5701
rect 11333 5661 11345 5695
rect 11379 5692 11391 5695
rect 12526 5692 12532 5704
rect 11379 5664 12532 5692
rect 11379 5661 11391 5664
rect 11333 5655 11391 5661
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 12618 5652 12624 5704
rect 12676 5692 12682 5704
rect 15378 5692 15384 5704
rect 12676 5664 15384 5692
rect 12676 5652 12682 5664
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 16025 5695 16083 5701
rect 16025 5661 16037 5695
rect 16071 5692 16083 5695
rect 16298 5692 16304 5704
rect 16071 5664 16304 5692
rect 16071 5661 16083 5664
rect 16025 5655 16083 5661
rect 16298 5652 16304 5664
rect 16356 5652 16362 5704
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5692 17187 5695
rect 20070 5692 20076 5704
rect 17175 5664 20076 5692
rect 17175 5661 17187 5664
rect 17129 5655 17187 5661
rect 20070 5652 20076 5664
rect 20128 5652 20134 5704
rect 23400 5692 23428 5723
rect 24854 5720 24860 5732
rect 24912 5720 24918 5772
rect 25222 5760 25228 5772
rect 25183 5732 25228 5760
rect 25222 5720 25228 5732
rect 25280 5720 25286 5772
rect 25314 5720 25320 5772
rect 25372 5760 25378 5772
rect 26804 5760 26832 5800
rect 26970 5760 26976 5772
rect 25372 5732 26832 5760
rect 26931 5732 26976 5760
rect 25372 5720 25378 5732
rect 26970 5720 26976 5732
rect 27028 5720 27034 5772
rect 27172 5769 27200 5800
rect 27157 5763 27215 5769
rect 27157 5729 27169 5763
rect 27203 5729 27215 5763
rect 27157 5723 27215 5729
rect 27246 5720 27252 5772
rect 27304 5720 27310 5772
rect 25041 5695 25099 5701
rect 25041 5692 25053 5695
rect 23400 5664 25053 5692
rect 25041 5661 25053 5664
rect 25087 5661 25099 5695
rect 27264 5692 27292 5720
rect 25041 5655 25099 5661
rect 26160 5664 27292 5692
rect 27356 5692 27384 5800
rect 27448 5800 27988 5828
rect 27448 5769 27476 5800
rect 27982 5788 27988 5800
rect 28040 5828 28046 5840
rect 28350 5828 28356 5840
rect 28040 5800 28356 5828
rect 28040 5788 28046 5800
rect 28350 5788 28356 5800
rect 28408 5788 28414 5840
rect 30190 5828 30196 5840
rect 28460 5800 30196 5828
rect 27433 5763 27491 5769
rect 27433 5729 27445 5763
rect 27479 5729 27491 5763
rect 27433 5723 27491 5729
rect 27522 5720 27528 5772
rect 27580 5760 27586 5772
rect 27617 5763 27675 5769
rect 27617 5760 27629 5763
rect 27580 5732 27629 5760
rect 27580 5720 27586 5732
rect 27617 5729 27629 5732
rect 27663 5729 27675 5763
rect 27617 5723 27675 5729
rect 27706 5720 27712 5772
rect 27764 5760 27770 5772
rect 27801 5763 27859 5769
rect 27801 5760 27813 5763
rect 27764 5732 27813 5760
rect 27764 5720 27770 5732
rect 27801 5729 27813 5732
rect 27847 5729 27859 5763
rect 27801 5723 27859 5729
rect 28460 5692 28488 5800
rect 30190 5788 30196 5800
rect 30248 5788 30254 5840
rect 32125 5831 32183 5837
rect 32125 5797 32137 5831
rect 32171 5828 32183 5831
rect 32398 5828 32404 5840
rect 32171 5800 32404 5828
rect 32171 5797 32183 5800
rect 32125 5791 32183 5797
rect 32398 5788 32404 5800
rect 32456 5828 32462 5840
rect 34606 5828 34612 5840
rect 32456 5800 34612 5828
rect 32456 5788 32462 5800
rect 34606 5788 34612 5800
rect 34664 5788 34670 5840
rect 34885 5831 34943 5837
rect 34885 5797 34897 5831
rect 34931 5828 34943 5831
rect 39114 5828 39120 5840
rect 34931 5800 39120 5828
rect 34931 5797 34943 5800
rect 34885 5791 34943 5797
rect 39114 5788 39120 5800
rect 39172 5788 39178 5840
rect 39482 5788 39488 5840
rect 39540 5828 39546 5840
rect 41340 5837 41368 5868
rect 42794 5856 42800 5868
rect 42852 5856 42858 5908
rect 42886 5856 42892 5908
rect 42944 5896 42950 5908
rect 42944 5868 47164 5896
rect 42944 5856 42950 5868
rect 41325 5831 41383 5837
rect 39540 5800 41092 5828
rect 39540 5788 39546 5800
rect 28905 5763 28963 5769
rect 28905 5729 28917 5763
rect 28951 5760 28963 5763
rect 30098 5760 30104 5772
rect 28951 5732 30104 5760
rect 28951 5729 28963 5732
rect 28905 5723 28963 5729
rect 30098 5720 30104 5732
rect 30156 5720 30162 5772
rect 30926 5720 30932 5772
rect 30984 5769 30990 5772
rect 30984 5763 31033 5769
rect 30984 5729 30987 5763
rect 31021 5729 31033 5763
rect 30984 5723 31033 5729
rect 30984 5720 30990 5723
rect 31110 5720 31116 5772
rect 31168 5760 31174 5772
rect 31205 5763 31263 5769
rect 31205 5760 31217 5763
rect 31168 5732 31217 5760
rect 31168 5720 31174 5732
rect 31205 5729 31217 5732
rect 31251 5729 31263 5763
rect 32306 5760 32312 5772
rect 32267 5732 32312 5760
rect 31205 5723 31263 5729
rect 32306 5720 32312 5732
rect 32364 5720 32370 5772
rect 32582 5720 32588 5772
rect 32640 5760 32646 5772
rect 34425 5763 34483 5769
rect 34425 5760 34437 5763
rect 32640 5732 34437 5760
rect 32640 5720 32646 5732
rect 34425 5729 34437 5732
rect 34471 5729 34483 5763
rect 34425 5723 34483 5729
rect 36449 5763 36507 5769
rect 36449 5729 36461 5763
rect 36495 5760 36507 5763
rect 37182 5760 37188 5772
rect 36495 5732 37188 5760
rect 36495 5729 36507 5732
rect 36449 5723 36507 5729
rect 37182 5720 37188 5732
rect 37240 5720 37246 5772
rect 37553 5763 37611 5769
rect 37553 5729 37565 5763
rect 37599 5760 37611 5763
rect 38105 5763 38163 5769
rect 38105 5760 38117 5763
rect 37599 5732 38117 5760
rect 37599 5729 37611 5732
rect 37553 5723 37611 5729
rect 38105 5729 38117 5732
rect 38151 5760 38163 5763
rect 38746 5760 38752 5772
rect 38151 5732 38752 5760
rect 38151 5729 38163 5732
rect 38105 5723 38163 5729
rect 38746 5720 38752 5732
rect 38804 5760 38810 5772
rect 39209 5763 39267 5769
rect 39209 5760 39221 5763
rect 38804 5732 39221 5760
rect 38804 5720 38810 5732
rect 39209 5729 39221 5732
rect 39255 5729 39267 5763
rect 39390 5760 39396 5772
rect 39351 5732 39396 5760
rect 39209 5723 39267 5729
rect 39390 5720 39396 5732
rect 39448 5720 39454 5772
rect 39761 5763 39819 5769
rect 39761 5729 39773 5763
rect 39807 5760 39819 5763
rect 40773 5763 40831 5769
rect 40773 5760 40785 5763
rect 39807 5732 40785 5760
rect 39807 5729 39819 5732
rect 39761 5723 39819 5729
rect 40773 5729 40785 5732
rect 40819 5729 40831 5763
rect 40773 5723 40831 5729
rect 40862 5720 40868 5772
rect 40920 5760 40926 5772
rect 41064 5760 41092 5800
rect 41325 5797 41337 5831
rect 41371 5797 41383 5831
rect 44634 5828 44640 5840
rect 41325 5791 41383 5797
rect 42076 5800 44640 5828
rect 42076 5760 42104 5800
rect 44634 5788 44640 5800
rect 44692 5788 44698 5840
rect 47029 5831 47087 5837
rect 47029 5828 47041 5831
rect 45388 5800 47041 5828
rect 40920 5732 40965 5760
rect 41064 5732 42104 5760
rect 42153 5763 42211 5769
rect 40920 5720 40926 5732
rect 42153 5729 42165 5763
rect 42199 5760 42211 5763
rect 42334 5760 42340 5772
rect 42199 5732 42340 5760
rect 42199 5729 42211 5732
rect 42153 5723 42211 5729
rect 42334 5720 42340 5732
rect 42392 5720 42398 5772
rect 43717 5763 43775 5769
rect 43717 5729 43729 5763
rect 43763 5760 43775 5763
rect 43809 5763 43867 5769
rect 43809 5760 43821 5763
rect 43763 5732 43821 5760
rect 43763 5729 43775 5732
rect 43717 5723 43775 5729
rect 43809 5729 43821 5732
rect 43855 5729 43867 5763
rect 43809 5723 43867 5729
rect 44082 5720 44088 5772
rect 44140 5760 44146 5772
rect 44177 5763 44235 5769
rect 44177 5760 44189 5763
rect 44140 5732 44189 5760
rect 44140 5720 44146 5732
rect 44177 5729 44189 5732
rect 44223 5729 44235 5763
rect 44450 5760 44456 5772
rect 44411 5732 44456 5760
rect 44177 5723 44235 5729
rect 44450 5720 44456 5732
rect 44508 5720 44514 5772
rect 45388 5769 45416 5800
rect 47029 5797 47041 5800
rect 47075 5797 47087 5831
rect 47136 5828 47164 5868
rect 47210 5856 47216 5908
rect 47268 5896 47274 5908
rect 48866 5896 48872 5908
rect 47268 5868 48872 5896
rect 47268 5856 47274 5868
rect 48866 5856 48872 5868
rect 48924 5856 48930 5908
rect 49418 5896 49424 5908
rect 49379 5868 49424 5896
rect 49418 5856 49424 5868
rect 49476 5856 49482 5908
rect 49528 5868 50016 5896
rect 49528 5828 49556 5868
rect 47136 5800 49556 5828
rect 49605 5831 49663 5837
rect 47029 5791 47087 5797
rect 49605 5797 49617 5831
rect 49651 5828 49663 5831
rect 49878 5828 49884 5840
rect 49651 5800 49884 5828
rect 49651 5797 49663 5800
rect 49605 5791 49663 5797
rect 49878 5788 49884 5800
rect 49936 5788 49942 5840
rect 49988 5837 50016 5868
rect 50246 5856 50252 5908
rect 50304 5896 50310 5908
rect 50522 5896 50528 5908
rect 50304 5868 50528 5896
rect 50304 5856 50310 5868
rect 50522 5856 50528 5868
rect 50580 5896 50586 5908
rect 52454 5896 52460 5908
rect 50580 5868 52460 5896
rect 50580 5856 50586 5868
rect 52454 5856 52460 5868
rect 52512 5856 52518 5908
rect 52822 5896 52828 5908
rect 52564 5868 52828 5896
rect 49973 5831 50031 5837
rect 49973 5797 49985 5831
rect 50019 5797 50031 5831
rect 49973 5791 50031 5797
rect 50614 5788 50620 5840
rect 50672 5828 50678 5840
rect 51534 5828 51540 5840
rect 50672 5800 51540 5828
rect 50672 5788 50678 5800
rect 51534 5788 51540 5800
rect 51592 5788 51598 5840
rect 52564 5828 52592 5868
rect 52822 5856 52828 5868
rect 52880 5896 52886 5908
rect 53101 5899 53159 5905
rect 53101 5896 53113 5899
rect 52880 5868 53113 5896
rect 52880 5856 52886 5868
rect 53101 5865 53113 5868
rect 53147 5865 53159 5899
rect 56502 5896 56508 5908
rect 53101 5859 53159 5865
rect 53208 5868 56508 5896
rect 51736 5800 52592 5828
rect 52917 5831 52975 5837
rect 45378 5763 45436 5769
rect 45378 5729 45390 5763
rect 45424 5729 45436 5763
rect 45646 5760 45652 5772
rect 45607 5732 45652 5760
rect 45378 5723 45436 5729
rect 45646 5720 45652 5732
rect 45704 5720 45710 5772
rect 47857 5763 47915 5769
rect 46032 5732 47808 5760
rect 27356 5664 28488 5692
rect 28813 5695 28871 5701
rect 6914 5624 6920 5636
rect 6875 5596 6920 5624
rect 6914 5584 6920 5596
rect 6972 5584 6978 5636
rect 8021 5627 8079 5633
rect 8021 5593 8033 5627
rect 8067 5624 8079 5627
rect 10962 5624 10968 5636
rect 8067 5596 10968 5624
rect 8067 5593 8079 5596
rect 8021 5587 8079 5593
rect 10962 5584 10968 5596
rect 11020 5584 11026 5636
rect 15286 5624 15292 5636
rect 11992 5596 15292 5624
rect 11992 5556 12020 5596
rect 15286 5584 15292 5596
rect 15344 5584 15350 5636
rect 22370 5584 22376 5636
rect 22428 5624 22434 5636
rect 26160 5624 26188 5664
rect 28813 5661 28825 5695
rect 28859 5692 28871 5695
rect 29270 5692 29276 5704
rect 28859 5664 29276 5692
rect 28859 5661 28871 5664
rect 28813 5655 28871 5661
rect 29270 5652 29276 5664
rect 29328 5652 29334 5704
rect 30190 5692 30196 5704
rect 30151 5664 30196 5692
rect 30190 5652 30196 5664
rect 30248 5652 30254 5704
rect 30466 5652 30472 5704
rect 30524 5692 30530 5704
rect 30745 5695 30803 5701
rect 30745 5692 30757 5695
rect 30524 5664 30757 5692
rect 30524 5652 30530 5664
rect 30745 5661 30757 5664
rect 30791 5661 30803 5695
rect 32674 5692 32680 5704
rect 32635 5664 32680 5692
rect 30745 5655 30803 5661
rect 32674 5652 32680 5664
rect 32732 5652 32738 5704
rect 33226 5652 33232 5704
rect 33284 5692 33290 5704
rect 34054 5692 34060 5704
rect 33284 5664 34060 5692
rect 33284 5652 33290 5664
rect 34054 5652 34060 5664
rect 34112 5652 34118 5704
rect 34330 5692 34336 5704
rect 34291 5664 34336 5692
rect 34330 5652 34336 5664
rect 34388 5652 34394 5704
rect 45186 5692 45192 5704
rect 34440 5664 45192 5692
rect 22428 5596 26188 5624
rect 22428 5584 22434 5596
rect 26418 5584 26424 5636
rect 26476 5624 26482 5636
rect 27706 5624 27712 5636
rect 26476 5596 27712 5624
rect 26476 5584 26482 5596
rect 27706 5584 27712 5596
rect 27764 5624 27770 5636
rect 27764 5596 31800 5624
rect 27764 5584 27770 5596
rect 6564 5528 12020 5556
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 13722 5556 13728 5568
rect 12492 5528 12537 5556
rect 13683 5528 13728 5556
rect 12492 5516 12498 5528
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 15470 5516 15476 5568
rect 15528 5556 15534 5568
rect 17494 5556 17500 5568
rect 15528 5528 17500 5556
rect 15528 5516 15534 5528
rect 17494 5516 17500 5528
rect 17552 5516 17558 5568
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 18233 5559 18291 5565
rect 18233 5556 18245 5559
rect 18012 5528 18245 5556
rect 18012 5516 18018 5528
rect 18233 5525 18245 5528
rect 18279 5525 18291 5559
rect 18233 5519 18291 5525
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 19613 5559 19671 5565
rect 19613 5556 19625 5559
rect 19392 5528 19625 5556
rect 19392 5516 19398 5528
rect 19613 5525 19625 5528
rect 19659 5525 19671 5559
rect 23106 5556 23112 5568
rect 23067 5528 23112 5556
rect 19613 5519 19671 5525
rect 23106 5516 23112 5528
rect 23164 5516 23170 5568
rect 23566 5556 23572 5568
rect 23527 5528 23572 5556
rect 23566 5516 23572 5528
rect 23624 5516 23630 5568
rect 23842 5516 23848 5568
rect 23900 5556 23906 5568
rect 28810 5556 28816 5568
rect 23900 5528 28816 5556
rect 23900 5516 23906 5528
rect 28810 5516 28816 5528
rect 28868 5516 28874 5568
rect 29086 5556 29092 5568
rect 29047 5528 29092 5556
rect 29086 5516 29092 5528
rect 29144 5516 29150 5568
rect 31772 5556 31800 5596
rect 31846 5584 31852 5636
rect 31904 5624 31910 5636
rect 34440 5624 34468 5664
rect 45186 5652 45192 5664
rect 45244 5652 45250 5704
rect 45462 5692 45468 5704
rect 45423 5664 45468 5692
rect 45462 5652 45468 5664
rect 45520 5652 45526 5704
rect 46032 5692 46060 5732
rect 45572 5664 46060 5692
rect 46109 5695 46167 5701
rect 31904 5596 34468 5624
rect 31904 5584 31910 5596
rect 34514 5584 34520 5636
rect 34572 5624 34578 5636
rect 36170 5624 36176 5636
rect 34572 5596 36176 5624
rect 34572 5584 34578 5596
rect 36170 5584 36176 5596
rect 36228 5584 36234 5636
rect 36354 5584 36360 5636
rect 36412 5624 36418 5636
rect 45572 5624 45600 5664
rect 46109 5661 46121 5695
rect 46155 5692 46167 5695
rect 46382 5692 46388 5704
rect 46155 5664 46388 5692
rect 46155 5661 46167 5664
rect 46109 5655 46167 5661
rect 46382 5652 46388 5664
rect 46440 5652 46446 5704
rect 47581 5695 47639 5701
rect 47581 5661 47593 5695
rect 47627 5661 47639 5695
rect 47780 5692 47808 5732
rect 47857 5729 47869 5763
rect 47903 5760 47915 5763
rect 49513 5763 49571 5769
rect 47903 5732 49372 5760
rect 47903 5729 47915 5732
rect 47857 5723 47915 5729
rect 48038 5692 48044 5704
rect 47780 5664 48044 5692
rect 47581 5655 47639 5661
rect 36412 5596 45600 5624
rect 36412 5584 36418 5596
rect 45646 5584 45652 5636
rect 45704 5624 45710 5636
rect 47210 5624 47216 5636
rect 45704 5596 47216 5624
rect 45704 5584 45710 5596
rect 47210 5584 47216 5596
rect 47268 5584 47274 5636
rect 47596 5624 47624 5655
rect 48038 5652 48044 5664
rect 48096 5652 48102 5704
rect 48130 5652 48136 5704
rect 48188 5692 48194 5704
rect 49234 5692 49240 5704
rect 48188 5664 49240 5692
rect 48188 5652 48194 5664
rect 49234 5652 49240 5664
rect 49292 5652 49298 5704
rect 49344 5692 49372 5732
rect 49513 5729 49525 5763
rect 49559 5760 49571 5763
rect 50430 5760 50436 5772
rect 49559 5732 50436 5760
rect 49559 5729 49571 5732
rect 49513 5723 49571 5729
rect 50430 5720 50436 5732
rect 50488 5760 50494 5772
rect 51258 5760 51264 5772
rect 50488 5732 51264 5760
rect 50488 5720 50494 5732
rect 51258 5720 51264 5732
rect 51316 5720 51322 5772
rect 51736 5769 51764 5800
rect 52917 5797 52929 5831
rect 52963 5828 52975 5831
rect 53208 5828 53236 5868
rect 56502 5856 56508 5868
rect 56560 5856 56566 5908
rect 57514 5856 57520 5908
rect 57572 5896 57578 5908
rect 57572 5868 60136 5896
rect 57572 5856 57578 5868
rect 52963 5800 53236 5828
rect 53285 5831 53343 5837
rect 52963 5797 52975 5800
rect 52917 5791 52975 5797
rect 53285 5797 53297 5831
rect 53331 5828 53343 5831
rect 53466 5828 53472 5840
rect 53331 5800 53472 5828
rect 53331 5797 53343 5800
rect 53285 5791 53343 5797
rect 53466 5788 53472 5800
rect 53524 5788 53530 5840
rect 55309 5831 55367 5837
rect 55309 5797 55321 5831
rect 55355 5828 55367 5831
rect 55398 5828 55404 5840
rect 55355 5800 55404 5828
rect 55355 5797 55367 5800
rect 55309 5791 55367 5797
rect 55398 5788 55404 5800
rect 55456 5828 55462 5840
rect 58437 5831 58495 5837
rect 55456 5800 57928 5828
rect 55456 5788 55462 5800
rect 51721 5763 51779 5769
rect 51721 5729 51733 5763
rect 51767 5729 51779 5763
rect 51721 5723 51779 5729
rect 49786 5692 49792 5704
rect 49344 5664 49792 5692
rect 49786 5652 49792 5664
rect 49844 5652 49850 5704
rect 47670 5624 47676 5636
rect 47583 5596 47676 5624
rect 47670 5584 47676 5596
rect 47728 5624 47734 5636
rect 51736 5624 51764 5723
rect 52086 5720 52092 5772
rect 52144 5760 52150 5772
rect 53193 5763 53251 5769
rect 52144 5732 53144 5760
rect 52144 5720 52150 5732
rect 53116 5692 53144 5732
rect 53193 5729 53205 5763
rect 53239 5760 53251 5763
rect 53374 5760 53380 5772
rect 53239 5732 53380 5760
rect 53239 5729 53251 5732
rect 53193 5723 53251 5729
rect 53374 5720 53380 5732
rect 53432 5720 53438 5772
rect 56137 5763 56195 5769
rect 56137 5760 56149 5763
rect 53484 5732 56149 5760
rect 53484 5692 53512 5732
rect 56137 5729 56149 5732
rect 56183 5760 56195 5763
rect 57149 5763 57207 5769
rect 57149 5760 57161 5763
rect 56183 5732 57161 5760
rect 56183 5729 56195 5732
rect 56137 5723 56195 5729
rect 57149 5729 57161 5732
rect 57195 5729 57207 5763
rect 57149 5723 57207 5729
rect 57333 5763 57391 5769
rect 57333 5729 57345 5763
rect 57379 5729 57391 5763
rect 57790 5760 57796 5772
rect 57751 5732 57796 5760
rect 57333 5723 57391 5729
rect 53116 5664 53512 5692
rect 53653 5695 53711 5701
rect 53653 5661 53665 5695
rect 53699 5661 53711 5695
rect 53653 5655 53711 5661
rect 52086 5624 52092 5636
rect 47728 5596 51764 5624
rect 51828 5596 52092 5624
rect 47728 5584 47734 5596
rect 36262 5556 36268 5568
rect 31772 5528 36268 5556
rect 36262 5516 36268 5528
rect 36320 5516 36326 5568
rect 36633 5559 36691 5565
rect 36633 5525 36645 5559
rect 36679 5556 36691 5559
rect 37274 5556 37280 5568
rect 36679 5528 37280 5556
rect 36679 5525 36691 5528
rect 36633 5519 36691 5525
rect 37274 5516 37280 5528
rect 37332 5516 37338 5568
rect 40586 5556 40592 5568
rect 40547 5528 40592 5556
rect 40586 5516 40592 5528
rect 40644 5516 40650 5568
rect 42058 5516 42064 5568
rect 42116 5556 42122 5568
rect 42337 5559 42395 5565
rect 42337 5556 42349 5559
rect 42116 5528 42349 5556
rect 42116 5516 42122 5528
rect 42337 5525 42349 5528
rect 42383 5556 42395 5559
rect 42426 5556 42432 5568
rect 42383 5528 42432 5556
rect 42383 5525 42395 5528
rect 42337 5519 42395 5525
rect 42426 5516 42432 5528
rect 42484 5516 42490 5568
rect 51828 5565 51856 5596
rect 52086 5584 52092 5596
rect 52144 5584 52150 5636
rect 52362 5584 52368 5636
rect 52420 5624 52426 5636
rect 53668 5624 53696 5655
rect 54754 5652 54760 5704
rect 54812 5692 54818 5704
rect 55861 5695 55919 5701
rect 55861 5692 55873 5695
rect 54812 5664 55873 5692
rect 54812 5652 54818 5664
rect 55861 5661 55873 5664
rect 55907 5661 55919 5695
rect 55861 5655 55919 5661
rect 56226 5652 56232 5704
rect 56284 5692 56290 5704
rect 56321 5695 56379 5701
rect 56321 5692 56333 5695
rect 56284 5664 56333 5692
rect 56284 5652 56290 5664
rect 56321 5661 56333 5664
rect 56367 5692 56379 5695
rect 57348 5692 57376 5723
rect 57790 5720 57796 5732
rect 57848 5720 57854 5772
rect 57900 5769 57928 5800
rect 58437 5797 58449 5831
rect 58483 5828 58495 5831
rect 59170 5828 59176 5840
rect 58483 5800 59176 5828
rect 58483 5797 58495 5800
rect 58437 5791 58495 5797
rect 59170 5788 59176 5800
rect 59228 5788 59234 5840
rect 57885 5763 57943 5769
rect 57885 5729 57897 5763
rect 57931 5729 57943 5763
rect 60108 5760 60136 5868
rect 60185 5763 60243 5769
rect 60185 5760 60197 5763
rect 60108 5732 60197 5760
rect 57885 5723 57943 5729
rect 60185 5729 60197 5732
rect 60231 5729 60243 5763
rect 60185 5723 60243 5729
rect 60277 5763 60335 5769
rect 60277 5729 60289 5763
rect 60323 5729 60335 5763
rect 60277 5723 60335 5729
rect 57514 5692 57520 5704
rect 56367 5664 57520 5692
rect 56367 5661 56379 5664
rect 56321 5655 56379 5661
rect 57514 5652 57520 5664
rect 57572 5652 57578 5704
rect 52420 5596 53696 5624
rect 52420 5584 52426 5596
rect 53834 5584 53840 5636
rect 53892 5624 53898 5636
rect 54386 5624 54392 5636
rect 53892 5596 54392 5624
rect 53892 5584 53898 5596
rect 54386 5584 54392 5596
rect 54444 5624 54450 5636
rect 54444 5596 56456 5624
rect 54444 5584 54450 5596
rect 43717 5559 43775 5565
rect 43717 5525 43729 5559
rect 43763 5556 43775 5559
rect 51813 5559 51871 5565
rect 51813 5556 51825 5559
rect 43763 5528 51825 5556
rect 43763 5525 43775 5528
rect 43717 5519 43775 5525
rect 51813 5525 51825 5528
rect 51859 5525 51871 5559
rect 51813 5519 51871 5525
rect 52270 5516 52276 5568
rect 52328 5556 52334 5568
rect 56318 5556 56324 5568
rect 52328 5528 56324 5556
rect 52328 5516 52334 5528
rect 56318 5516 56324 5528
rect 56376 5516 56382 5568
rect 56428 5556 56456 5596
rect 57698 5584 57704 5636
rect 57756 5624 57762 5636
rect 60292 5624 60320 5723
rect 57756 5596 60320 5624
rect 57756 5584 57762 5596
rect 58342 5556 58348 5568
rect 56428 5528 58348 5556
rect 58342 5516 58348 5528
rect 58400 5556 58406 5568
rect 58618 5556 58624 5568
rect 58400 5528 58624 5556
rect 58400 5516 58406 5528
rect 58618 5516 58624 5528
rect 58676 5516 58682 5568
rect 58802 5516 58808 5568
rect 58860 5556 58866 5568
rect 60461 5559 60519 5565
rect 60461 5556 60473 5559
rect 58860 5528 60473 5556
rect 58860 5516 58866 5528
rect 60461 5525 60473 5528
rect 60507 5525 60519 5559
rect 60461 5519 60519 5525
rect 1104 5466 62192 5488
rect 1104 5414 11163 5466
rect 11215 5414 11227 5466
rect 11279 5414 11291 5466
rect 11343 5414 11355 5466
rect 11407 5414 31526 5466
rect 31578 5414 31590 5466
rect 31642 5414 31654 5466
rect 31706 5414 31718 5466
rect 31770 5414 51888 5466
rect 51940 5414 51952 5466
rect 52004 5414 52016 5466
rect 52068 5414 52080 5466
rect 52132 5414 62192 5466
rect 1104 5392 62192 5414
rect 2958 5312 2964 5364
rect 3016 5352 3022 5364
rect 3053 5355 3111 5361
rect 3053 5352 3065 5355
rect 3016 5324 3065 5352
rect 3016 5312 3022 5324
rect 3053 5321 3065 5324
rect 3099 5321 3111 5355
rect 3053 5315 3111 5321
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 6362 5352 6368 5364
rect 5767 5324 6368 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 7101 5355 7159 5361
rect 7101 5352 7113 5355
rect 7064 5324 7113 5352
rect 7064 5312 7070 5324
rect 7101 5321 7113 5324
rect 7147 5321 7159 5355
rect 12526 5352 12532 5364
rect 12487 5324 12532 5352
rect 7101 5315 7159 5321
rect 12526 5312 12532 5324
rect 12584 5312 12590 5364
rect 14918 5352 14924 5364
rect 13096 5324 14924 5352
rect 10597 5287 10655 5293
rect 7484 5256 10456 5284
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5216 2835 5219
rect 7484 5216 7512 5256
rect 2823 5188 7512 5216
rect 7561 5219 7619 5225
rect 2823 5185 2835 5188
rect 2777 5179 2835 5185
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 8386 5216 8392 5228
rect 7607 5188 8392 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 10428 5216 10456 5256
rect 10597 5253 10609 5287
rect 10643 5284 10655 5287
rect 13096 5284 13124 5324
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 16666 5312 16672 5364
rect 16724 5352 16730 5364
rect 17954 5352 17960 5364
rect 16724 5324 17960 5352
rect 16724 5312 16730 5324
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 18049 5355 18107 5361
rect 18049 5321 18061 5355
rect 18095 5352 18107 5355
rect 20898 5352 20904 5364
rect 18095 5324 20904 5352
rect 18095 5321 18107 5324
rect 18049 5315 18107 5321
rect 20898 5312 20904 5324
rect 20956 5352 20962 5364
rect 23106 5352 23112 5364
rect 20956 5324 23112 5352
rect 20956 5312 20962 5324
rect 23106 5312 23112 5324
rect 23164 5312 23170 5364
rect 25498 5312 25504 5364
rect 25556 5352 25562 5364
rect 36722 5352 36728 5364
rect 25556 5324 36728 5352
rect 25556 5312 25562 5324
rect 36722 5312 36728 5324
rect 36780 5352 36786 5364
rect 38010 5352 38016 5364
rect 36780 5324 38016 5352
rect 36780 5312 36786 5324
rect 38010 5312 38016 5324
rect 38068 5312 38074 5364
rect 40773 5355 40831 5361
rect 40773 5321 40785 5355
rect 40819 5352 40831 5355
rect 40862 5352 40868 5364
rect 40819 5324 40868 5352
rect 40819 5321 40831 5324
rect 40773 5315 40831 5321
rect 40862 5312 40868 5324
rect 40920 5312 40926 5364
rect 40954 5312 40960 5364
rect 41012 5352 41018 5364
rect 51442 5352 51448 5364
rect 41012 5324 43484 5352
rect 41012 5312 41018 5324
rect 23566 5284 23572 5296
rect 10643 5256 13124 5284
rect 13188 5256 23572 5284
rect 10643 5253 10655 5256
rect 10597 5247 10655 5253
rect 11054 5216 11060 5228
rect 10428 5188 11060 5216
rect 11054 5176 11060 5188
rect 11112 5176 11118 5228
rect 11333 5219 11391 5225
rect 11333 5185 11345 5219
rect 11379 5216 11391 5219
rect 12250 5216 12256 5228
rect 11379 5188 12256 5216
rect 11379 5185 11391 5188
rect 11333 5179 11391 5185
rect 12250 5176 12256 5188
rect 12308 5176 12314 5228
rect 13188 5225 13216 5256
rect 23566 5244 23572 5256
rect 23624 5244 23630 5296
rect 24121 5287 24179 5293
rect 24121 5253 24133 5287
rect 24167 5253 24179 5287
rect 26878 5284 26884 5296
rect 26839 5256 26884 5284
rect 24121 5247 24179 5253
rect 13173 5219 13231 5225
rect 13173 5185 13185 5219
rect 13219 5185 13231 5219
rect 13722 5216 13728 5228
rect 13173 5179 13231 5185
rect 13464 5188 13728 5216
rect 2866 5108 2872 5160
rect 2924 5157 2930 5160
rect 2924 5151 2947 5157
rect 2935 5117 2947 5151
rect 4154 5148 4160 5160
rect 4115 5120 4160 5148
rect 2924 5111 2947 5117
rect 2924 5108 2930 5111
rect 4154 5108 4160 5120
rect 4212 5108 4218 5160
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 5350 5148 5356 5160
rect 4479 5120 5356 5148
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 7469 5151 7527 5157
rect 7469 5148 7481 5151
rect 7340 5120 7481 5148
rect 7340 5108 7346 5120
rect 7469 5117 7481 5120
rect 7515 5117 7527 5151
rect 7834 5148 7840 5160
rect 7795 5120 7840 5148
rect 7469 5111 7527 5117
rect 7834 5108 7840 5120
rect 7892 5108 7898 5160
rect 8021 5151 8079 5157
rect 8021 5117 8033 5151
rect 8067 5148 8079 5151
rect 8202 5148 8208 5160
rect 8067 5120 8208 5148
rect 8067 5117 8079 5120
rect 8021 5111 8079 5117
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 8938 5108 8944 5160
rect 8996 5148 9002 5160
rect 9033 5151 9091 5157
rect 9033 5148 9045 5151
rect 8996 5120 9045 5148
rect 8996 5108 9002 5120
rect 9033 5117 9045 5120
rect 9079 5148 9091 5151
rect 9122 5148 9128 5160
rect 9079 5120 9128 5148
rect 9079 5117 9091 5120
rect 9033 5111 9091 5117
rect 9122 5108 9128 5120
rect 9180 5108 9186 5160
rect 10870 5148 10876 5160
rect 10831 5120 10876 5148
rect 10870 5108 10876 5120
rect 10928 5108 10934 5160
rect 13078 5148 13084 5160
rect 13039 5120 13084 5148
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13464 5157 13492 5188
rect 13722 5176 13728 5188
rect 13780 5176 13786 5228
rect 15286 5216 15292 5228
rect 15247 5188 15292 5216
rect 15286 5176 15292 5188
rect 15344 5176 15350 5228
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 18785 5219 18843 5225
rect 16163 5188 18460 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 13449 5151 13507 5157
rect 13449 5117 13461 5151
rect 13495 5117 13507 5151
rect 13449 5111 13507 5117
rect 13538 5108 13544 5160
rect 13596 5148 13602 5160
rect 14737 5151 14795 5157
rect 13596 5120 13641 5148
rect 13596 5108 13602 5120
rect 14737 5117 14749 5151
rect 14783 5117 14795 5151
rect 14737 5111 14795 5117
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5148 14887 5151
rect 15194 5148 15200 5160
rect 14875 5120 15200 5148
rect 14875 5117 14887 5120
rect 14829 5111 14887 5117
rect 5718 5040 5724 5092
rect 5776 5080 5782 5092
rect 8849 5083 8907 5089
rect 8849 5080 8861 5083
rect 5776 5052 8861 5080
rect 5776 5040 5782 5052
rect 8849 5049 8861 5052
rect 8895 5080 8907 5083
rect 10781 5083 10839 5089
rect 8895 5052 9260 5080
rect 8895 5049 8907 5052
rect 8849 5043 8907 5049
rect 7926 4972 7932 5024
rect 7984 5012 7990 5024
rect 9125 5015 9183 5021
rect 9125 5012 9137 5015
rect 7984 4984 9137 5012
rect 7984 4972 7990 4984
rect 9125 4981 9137 4984
rect 9171 4981 9183 5015
rect 9232 5012 9260 5052
rect 10781 5049 10793 5083
rect 10827 5080 10839 5083
rect 14090 5080 14096 5092
rect 10827 5052 14096 5080
rect 10827 5049 10839 5052
rect 10781 5043 10839 5049
rect 14090 5040 14096 5052
rect 14148 5040 14154 5092
rect 13722 5012 13728 5024
rect 9232 4984 13728 5012
rect 9125 4975 9183 4981
rect 13722 4972 13728 4984
rect 13780 4972 13786 5024
rect 14752 5012 14780 5111
rect 15194 5108 15200 5120
rect 15252 5108 15258 5160
rect 15304 5080 15332 5176
rect 15746 5108 15752 5160
rect 15804 5148 15810 5160
rect 16666 5148 16672 5160
rect 15804 5120 16672 5148
rect 15804 5108 15810 5120
rect 16666 5108 16672 5120
rect 16724 5108 16730 5160
rect 16945 5151 17003 5157
rect 16945 5117 16957 5151
rect 16991 5117 17003 5151
rect 16945 5111 17003 5117
rect 17129 5151 17187 5157
rect 17129 5117 17141 5151
rect 17175 5148 17187 5151
rect 17218 5148 17224 5160
rect 17175 5120 17224 5148
rect 17175 5117 17187 5120
rect 17129 5111 17187 5117
rect 16960 5080 16988 5111
rect 17218 5108 17224 5120
rect 17276 5108 17282 5160
rect 18325 5151 18383 5157
rect 18325 5117 18337 5151
rect 18371 5117 18383 5151
rect 18432 5148 18460 5188
rect 18785 5185 18797 5219
rect 18831 5216 18843 5219
rect 19705 5219 19763 5225
rect 19705 5216 19717 5219
rect 18831 5188 19717 5216
rect 18831 5185 18843 5188
rect 18785 5179 18843 5185
rect 19705 5185 19717 5188
rect 19751 5185 19763 5219
rect 20070 5216 20076 5228
rect 20031 5188 20076 5216
rect 19705 5179 19763 5185
rect 20070 5176 20076 5188
rect 20128 5176 20134 5228
rect 20622 5176 20628 5228
rect 20680 5216 20686 5228
rect 24136 5216 24164 5247
rect 26878 5244 26884 5256
rect 26936 5244 26942 5296
rect 26970 5244 26976 5296
rect 27028 5284 27034 5296
rect 28442 5284 28448 5296
rect 27028 5256 28448 5284
rect 27028 5244 27034 5256
rect 28442 5244 28448 5256
rect 28500 5284 28506 5296
rect 43456 5293 43484 5324
rect 45572 5324 51448 5352
rect 30469 5287 30527 5293
rect 30469 5284 30481 5287
rect 28500 5256 30481 5284
rect 28500 5244 28506 5256
rect 30469 5253 30481 5256
rect 30515 5253 30527 5287
rect 43441 5287 43499 5293
rect 30469 5247 30527 5253
rect 31772 5256 42472 5284
rect 20680 5188 24164 5216
rect 20680 5176 20686 5188
rect 24302 5176 24308 5228
rect 24360 5216 24366 5228
rect 31772 5216 31800 5256
rect 32674 5216 32680 5228
rect 24360 5188 31800 5216
rect 31864 5188 32680 5216
rect 24360 5176 24366 5188
rect 19613 5151 19671 5157
rect 19613 5148 19625 5151
rect 18432 5120 19625 5148
rect 18325 5111 18383 5117
rect 19613 5117 19625 5120
rect 19659 5117 19671 5151
rect 19886 5148 19892 5160
rect 19847 5120 19892 5148
rect 19613 5111 19671 5117
rect 18230 5080 18236 5092
rect 15304 5052 16988 5080
rect 18191 5052 18236 5080
rect 18230 5040 18236 5052
rect 18288 5040 18294 5092
rect 18340 5080 18368 5111
rect 19886 5108 19892 5120
rect 19944 5108 19950 5160
rect 19978 5108 19984 5160
rect 20036 5148 20042 5160
rect 21361 5151 21419 5157
rect 21361 5148 21373 5151
rect 20036 5120 21373 5148
rect 20036 5108 20042 5120
rect 21361 5117 21373 5120
rect 21407 5117 21419 5151
rect 24026 5148 24032 5160
rect 23987 5120 24032 5148
rect 21361 5111 21419 5117
rect 24026 5108 24032 5120
rect 24084 5108 24090 5160
rect 24489 5151 24547 5157
rect 24489 5117 24501 5151
rect 24535 5117 24547 5151
rect 24489 5111 24547 5117
rect 25225 5151 25283 5157
rect 25225 5117 25237 5151
rect 25271 5148 25283 5151
rect 25314 5148 25320 5160
rect 25271 5120 25320 5148
rect 25271 5117 25283 5120
rect 25225 5111 25283 5117
rect 21174 5080 21180 5092
rect 18340 5052 20208 5080
rect 21135 5052 21180 5080
rect 15562 5012 15568 5024
rect 14752 4984 15568 5012
rect 15562 4972 15568 4984
rect 15620 4972 15626 5024
rect 15654 4972 15660 5024
rect 15712 5012 15718 5024
rect 17862 5012 17868 5024
rect 15712 4984 17868 5012
rect 15712 4972 15718 4984
rect 17862 4972 17868 4984
rect 17920 4972 17926 5024
rect 20180 5012 20208 5052
rect 21174 5040 21180 5052
rect 21232 5040 21238 5092
rect 23658 5040 23664 5092
rect 23716 5080 23722 5092
rect 24504 5080 24532 5111
rect 25314 5108 25320 5120
rect 25372 5108 25378 5160
rect 25498 5148 25504 5160
rect 25459 5120 25504 5148
rect 25498 5108 25504 5120
rect 25556 5108 25562 5160
rect 25958 5148 25964 5160
rect 25919 5120 25964 5148
rect 25958 5108 25964 5120
rect 26016 5108 26022 5160
rect 26602 5108 26608 5160
rect 26660 5148 26666 5160
rect 26789 5151 26847 5157
rect 26789 5148 26801 5151
rect 26660 5120 26801 5148
rect 26660 5108 26666 5120
rect 26789 5117 26801 5120
rect 26835 5117 26847 5151
rect 26789 5111 26847 5117
rect 27341 5151 27399 5157
rect 27341 5117 27353 5151
rect 27387 5117 27399 5151
rect 27341 5111 27399 5117
rect 30285 5151 30343 5157
rect 30285 5117 30297 5151
rect 30331 5117 30343 5151
rect 30285 5111 30343 5117
rect 31573 5151 31631 5157
rect 31573 5117 31585 5151
rect 31619 5148 31631 5151
rect 31864 5148 31892 5188
rect 32674 5176 32680 5188
rect 32732 5176 32738 5228
rect 35897 5219 35955 5225
rect 35897 5185 35909 5219
rect 35943 5216 35955 5219
rect 40586 5216 40592 5228
rect 35943 5188 40592 5216
rect 35943 5185 35955 5188
rect 35897 5179 35955 5185
rect 40586 5176 40592 5188
rect 40644 5216 40650 5228
rect 40954 5216 40960 5228
rect 40644 5188 40960 5216
rect 40644 5176 40650 5188
rect 40954 5176 40960 5188
rect 41012 5176 41018 5228
rect 41598 5216 41604 5228
rect 41064 5188 41604 5216
rect 31619 5120 31892 5148
rect 31619 5117 31631 5120
rect 31573 5111 31631 5117
rect 27356 5080 27384 5111
rect 27706 5080 27712 5092
rect 23716 5052 27712 5080
rect 23716 5040 23722 5052
rect 27706 5040 27712 5052
rect 27764 5040 27770 5092
rect 30300 5080 30328 5111
rect 31938 5108 31944 5160
rect 31996 5148 32002 5160
rect 32214 5148 32220 5160
rect 31996 5120 32041 5148
rect 32175 5120 32220 5148
rect 31996 5108 32002 5120
rect 32214 5108 32220 5120
rect 32272 5108 32278 5160
rect 32306 5108 32312 5160
rect 32364 5148 32370 5160
rect 32490 5148 32496 5160
rect 32364 5120 32496 5148
rect 32364 5108 32370 5120
rect 32490 5108 32496 5120
rect 32548 5108 32554 5160
rect 33318 5148 33324 5160
rect 33279 5120 33324 5148
rect 33318 5108 33324 5120
rect 33376 5108 33382 5160
rect 34790 5108 34796 5160
rect 34848 5148 34854 5160
rect 34885 5151 34943 5157
rect 34885 5148 34897 5151
rect 34848 5120 34897 5148
rect 34848 5108 34854 5120
rect 34885 5117 34897 5120
rect 34931 5117 34943 5151
rect 36446 5148 36452 5160
rect 36407 5120 36452 5148
rect 34885 5111 34943 5117
rect 36446 5108 36452 5120
rect 36504 5108 36510 5160
rect 36538 5108 36544 5160
rect 36596 5148 36602 5160
rect 36722 5148 36728 5160
rect 36596 5120 36641 5148
rect 36683 5120 36728 5148
rect 36596 5108 36602 5120
rect 36722 5108 36728 5120
rect 36780 5108 36786 5160
rect 36906 5148 36912 5160
rect 36867 5120 36912 5148
rect 36906 5108 36912 5120
rect 36964 5148 36970 5160
rect 37090 5148 37096 5160
rect 36964 5120 37096 5148
rect 36964 5108 36970 5120
rect 37090 5108 37096 5120
rect 37148 5108 37154 5160
rect 37182 5108 37188 5160
rect 37240 5148 37246 5160
rect 37277 5151 37335 5157
rect 37277 5148 37289 5151
rect 37240 5120 37289 5148
rect 37240 5108 37246 5120
rect 37277 5117 37289 5120
rect 37323 5117 37335 5151
rect 39022 5148 39028 5160
rect 38983 5120 39028 5148
rect 37277 5111 37335 5117
rect 39022 5108 39028 5120
rect 39080 5108 39086 5160
rect 39114 5108 39120 5160
rect 39172 5148 39178 5160
rect 39209 5151 39267 5157
rect 39209 5148 39221 5151
rect 39172 5120 39221 5148
rect 39172 5108 39178 5120
rect 39209 5117 39221 5120
rect 39255 5148 39267 5151
rect 39482 5148 39488 5160
rect 39255 5120 39488 5148
rect 39255 5117 39267 5120
rect 39209 5111 39267 5117
rect 39482 5108 39488 5120
rect 39540 5108 39546 5160
rect 39577 5151 39635 5157
rect 39577 5117 39589 5151
rect 39623 5148 39635 5151
rect 39666 5148 39672 5160
rect 39623 5120 39672 5148
rect 39623 5117 39635 5120
rect 39577 5111 39635 5117
rect 39666 5108 39672 5120
rect 39724 5108 39730 5160
rect 40310 5108 40316 5160
rect 40368 5148 40374 5160
rect 40681 5151 40739 5157
rect 40681 5148 40693 5151
rect 40368 5120 40693 5148
rect 40368 5108 40374 5120
rect 40681 5117 40693 5120
rect 40727 5148 40739 5151
rect 41064 5148 41092 5188
rect 41598 5176 41604 5188
rect 41656 5176 41662 5228
rect 41414 5148 41420 5160
rect 40727 5120 41092 5148
rect 41375 5120 41420 5148
rect 40727 5117 40739 5120
rect 40681 5111 40739 5117
rect 41414 5108 41420 5120
rect 41472 5108 41478 5160
rect 42242 5148 42248 5160
rect 42203 5120 42248 5148
rect 42242 5108 42248 5120
rect 42300 5108 42306 5160
rect 32858 5080 32864 5092
rect 30300 5052 32864 5080
rect 32858 5040 32864 5052
rect 32916 5040 32922 5092
rect 38930 5080 38936 5092
rect 33336 5052 38936 5080
rect 21453 5015 21511 5021
rect 21453 5012 21465 5015
rect 20180 4984 21465 5012
rect 21453 4981 21465 4984
rect 21499 4981 21511 5015
rect 21453 4975 21511 4981
rect 25958 4972 25964 5024
rect 26016 5012 26022 5024
rect 28718 5012 28724 5024
rect 26016 4984 28724 5012
rect 26016 4972 26022 4984
rect 28718 4972 28724 4984
rect 28776 4972 28782 5024
rect 30558 4972 30564 5024
rect 30616 5012 30622 5024
rect 31481 5015 31539 5021
rect 31481 5012 31493 5015
rect 30616 4984 31493 5012
rect 30616 4972 30622 4984
rect 31481 4981 31493 4984
rect 31527 5012 31539 5015
rect 33336 5012 33364 5052
rect 38930 5040 38936 5052
rect 38988 5040 38994 5092
rect 31527 4984 33364 5012
rect 31527 4981 31539 4984
rect 31481 4975 31539 4981
rect 33410 4972 33416 5024
rect 33468 5012 33474 5024
rect 33505 5015 33563 5021
rect 33505 5012 33517 5015
rect 33468 4984 33517 5012
rect 33468 4972 33474 4984
rect 33505 4981 33517 4984
rect 33551 5012 33563 5015
rect 34238 5012 34244 5024
rect 33551 4984 34244 5012
rect 33551 4981 33563 4984
rect 33505 4975 33563 4981
rect 34238 4972 34244 4984
rect 34296 4972 34302 5024
rect 34882 4972 34888 5024
rect 34940 5012 34946 5024
rect 34977 5015 35035 5021
rect 34977 5012 34989 5015
rect 34940 4984 34989 5012
rect 34940 4972 34946 4984
rect 34977 4981 34989 4984
rect 35023 4981 35035 5015
rect 34977 4975 35035 4981
rect 36170 4972 36176 5024
rect 36228 5012 36234 5024
rect 36906 5012 36912 5024
rect 36228 4984 36912 5012
rect 36228 4972 36234 4984
rect 36906 4972 36912 4984
rect 36964 4972 36970 5024
rect 42444 5021 42472 5256
rect 43441 5253 43453 5287
rect 43487 5284 43499 5287
rect 45572 5284 45600 5324
rect 51442 5312 51448 5324
rect 51500 5312 51506 5364
rect 51534 5312 51540 5364
rect 51592 5352 51598 5364
rect 53006 5352 53012 5364
rect 51592 5324 53012 5352
rect 51592 5312 51598 5324
rect 53006 5312 53012 5324
rect 53064 5312 53070 5364
rect 54573 5355 54631 5361
rect 54573 5321 54585 5355
rect 54619 5352 54631 5355
rect 55306 5352 55312 5364
rect 54619 5324 55312 5352
rect 54619 5321 54631 5324
rect 54573 5315 54631 5321
rect 55306 5312 55312 5324
rect 55364 5312 55370 5364
rect 57514 5312 57520 5364
rect 57572 5352 57578 5364
rect 57609 5355 57667 5361
rect 57609 5352 57621 5355
rect 57572 5324 57621 5352
rect 57572 5312 57578 5324
rect 57609 5321 57621 5324
rect 57655 5321 57667 5355
rect 57609 5315 57667 5321
rect 47670 5284 47676 5296
rect 43487 5256 45600 5284
rect 47631 5256 47676 5284
rect 43487 5253 43499 5256
rect 43441 5247 43499 5253
rect 47670 5244 47676 5256
rect 47728 5244 47734 5296
rect 50062 5284 50068 5296
rect 50023 5256 50068 5284
rect 50062 5244 50068 5256
rect 50120 5244 50126 5296
rect 52825 5287 52883 5293
rect 52825 5253 52837 5287
rect 52871 5284 52883 5287
rect 53466 5284 53472 5296
rect 52871 5256 53472 5284
rect 52871 5253 52883 5256
rect 52825 5247 52883 5253
rect 53466 5244 53472 5256
rect 53524 5244 53530 5296
rect 44177 5219 44235 5225
rect 44177 5185 44189 5219
rect 44223 5216 44235 5219
rect 45462 5216 45468 5228
rect 44223 5188 45468 5216
rect 44223 5185 44235 5188
rect 44177 5179 44235 5185
rect 45462 5176 45468 5188
rect 45520 5176 45526 5228
rect 46382 5216 46388 5228
rect 46343 5188 46388 5216
rect 46382 5176 46388 5188
rect 46440 5176 46446 5228
rect 46492 5188 50660 5216
rect 43714 5148 43720 5160
rect 43675 5120 43720 5148
rect 43714 5108 43720 5120
rect 43772 5108 43778 5160
rect 46106 5148 46112 5160
rect 46067 5120 46112 5148
rect 46106 5108 46112 5120
rect 46164 5108 46170 5160
rect 46198 5108 46204 5160
rect 46256 5148 46262 5160
rect 46492 5148 46520 5188
rect 46256 5120 46520 5148
rect 49421 5151 49479 5157
rect 46256 5108 46262 5120
rect 49421 5117 49433 5151
rect 49467 5148 49479 5151
rect 49602 5148 49608 5160
rect 49467 5120 49608 5148
rect 49467 5117 49479 5120
rect 49421 5111 49479 5117
rect 49602 5108 49608 5120
rect 49660 5108 49666 5160
rect 49786 5148 49792 5160
rect 49747 5120 49792 5148
rect 49786 5108 49792 5120
rect 49844 5108 49850 5160
rect 50065 5151 50123 5157
rect 50065 5117 50077 5151
rect 50111 5117 50123 5151
rect 50065 5111 50123 5117
rect 43625 5083 43683 5089
rect 43625 5049 43637 5083
rect 43671 5080 43683 5083
rect 44174 5080 44180 5092
rect 43671 5052 44180 5080
rect 43671 5049 43683 5052
rect 43625 5043 43683 5049
rect 44174 5040 44180 5052
rect 44232 5040 44238 5092
rect 42429 5015 42487 5021
rect 42429 4981 42441 5015
rect 42475 5012 42487 5015
rect 46216 5012 46244 5108
rect 47946 5040 47952 5092
rect 48004 5080 48010 5092
rect 50080 5080 50108 5111
rect 50430 5080 50436 5092
rect 48004 5052 50436 5080
rect 48004 5040 48010 5052
rect 50430 5040 50436 5052
rect 50488 5040 50494 5092
rect 42475 4984 46244 5012
rect 42475 4981 42487 4984
rect 42429 4975 42487 4981
rect 49970 4972 49976 5024
rect 50028 5012 50034 5024
rect 50522 5012 50528 5024
rect 50028 4984 50528 5012
rect 50028 4972 50034 4984
rect 50522 4972 50528 4984
rect 50580 4972 50586 5024
rect 50632 5012 50660 5188
rect 50798 5176 50804 5228
rect 50856 5216 50862 5228
rect 52917 5219 52975 5225
rect 52917 5216 52929 5219
rect 50856 5188 52929 5216
rect 50856 5176 50862 5188
rect 52917 5185 52929 5188
rect 52963 5216 52975 5219
rect 53374 5216 53380 5228
rect 52963 5188 53380 5216
rect 52963 5185 52975 5188
rect 52917 5179 52975 5185
rect 53374 5176 53380 5188
rect 53432 5176 53438 5228
rect 53484 5216 53512 5244
rect 57974 5216 57980 5228
rect 53484 5188 57980 5216
rect 52696 5151 52754 5157
rect 52696 5117 52708 5151
rect 52742 5148 52754 5151
rect 53742 5148 53748 5160
rect 52742 5120 53748 5148
rect 52742 5117 52754 5120
rect 52696 5111 52754 5117
rect 53742 5108 53748 5120
rect 53800 5108 53806 5160
rect 54573 5151 54631 5157
rect 54573 5117 54585 5151
rect 54619 5148 54631 5151
rect 54665 5151 54723 5157
rect 54665 5148 54677 5151
rect 54619 5120 54677 5148
rect 54619 5117 54631 5120
rect 54573 5111 54631 5117
rect 54665 5117 54677 5120
rect 54711 5117 54723 5151
rect 54665 5111 54723 5117
rect 54757 5151 54815 5157
rect 54757 5117 54769 5151
rect 54803 5148 54815 5151
rect 54846 5148 54852 5160
rect 54803 5120 54852 5148
rect 54803 5117 54815 5120
rect 54757 5111 54815 5117
rect 50706 5040 50712 5092
rect 50764 5080 50770 5092
rect 52549 5083 52607 5089
rect 52549 5080 52561 5083
rect 50764 5052 52561 5080
rect 50764 5040 50770 5052
rect 52549 5049 52561 5052
rect 52595 5049 52607 5083
rect 54772 5080 54800 5111
rect 54846 5108 54852 5120
rect 54904 5108 54910 5160
rect 54956 5157 54984 5188
rect 57974 5176 57980 5188
rect 58032 5176 58038 5228
rect 58066 5176 58072 5228
rect 58124 5216 58130 5228
rect 58805 5219 58863 5225
rect 58805 5216 58817 5219
rect 58124 5188 58817 5216
rect 58124 5176 58130 5188
rect 58805 5185 58817 5188
rect 58851 5185 58863 5219
rect 58805 5179 58863 5185
rect 54941 5151 54999 5157
rect 54941 5117 54953 5151
rect 54987 5117 54999 5151
rect 54941 5111 54999 5117
rect 56502 5108 56508 5160
rect 56560 5148 56566 5160
rect 57425 5151 57483 5157
rect 57425 5148 57437 5151
rect 56560 5120 57437 5148
rect 56560 5108 56566 5120
rect 57425 5117 57437 5120
rect 57471 5117 57483 5151
rect 57425 5111 57483 5117
rect 55398 5080 55404 5092
rect 52549 5043 52607 5049
rect 54680 5052 54800 5080
rect 55359 5052 55404 5080
rect 54680 5012 54708 5052
rect 55398 5040 55404 5052
rect 55456 5040 55462 5092
rect 50632 4984 54708 5012
rect 57440 5012 57468 5111
rect 58434 5108 58440 5160
rect 58492 5148 58498 5160
rect 58529 5151 58587 5157
rect 58529 5148 58541 5151
rect 58492 5120 58541 5148
rect 58492 5108 58498 5120
rect 58529 5117 58541 5120
rect 58575 5117 58587 5151
rect 58529 5111 58587 5117
rect 59909 5015 59967 5021
rect 59909 5012 59921 5015
rect 57440 4984 59921 5012
rect 59909 4981 59921 4984
rect 59955 4981 59967 5015
rect 59909 4975 59967 4981
rect 1104 4922 62192 4944
rect 1104 4870 21344 4922
rect 21396 4870 21408 4922
rect 21460 4870 21472 4922
rect 21524 4870 21536 4922
rect 21588 4870 41707 4922
rect 41759 4870 41771 4922
rect 41823 4870 41835 4922
rect 41887 4870 41899 4922
rect 41951 4870 62192 4922
rect 1104 4848 62192 4870
rect 6362 4768 6368 4820
rect 6420 4808 6426 4820
rect 11609 4811 11667 4817
rect 11609 4808 11621 4811
rect 6420 4780 11621 4808
rect 6420 4768 6426 4780
rect 11609 4777 11621 4780
rect 11655 4777 11667 4811
rect 11609 4771 11667 4777
rect 12345 4811 12403 4817
rect 12345 4777 12357 4811
rect 12391 4808 12403 4811
rect 15194 4808 15200 4820
rect 12391 4780 15200 4808
rect 12391 4777 12403 4780
rect 12345 4771 12403 4777
rect 15194 4768 15200 4780
rect 15252 4808 15258 4820
rect 15252 4780 15332 4808
rect 15252 4768 15258 4780
rect 3145 4743 3203 4749
rect 3145 4709 3157 4743
rect 3191 4740 3203 4743
rect 3234 4740 3240 4752
rect 3191 4712 3240 4740
rect 3191 4709 3203 4712
rect 3145 4703 3203 4709
rect 3234 4700 3240 4712
rect 3292 4700 3298 4752
rect 5350 4740 5356 4752
rect 5311 4712 5356 4740
rect 5350 4700 5356 4712
rect 5408 4700 5414 4752
rect 8386 4740 8392 4752
rect 7300 4712 8392 4740
rect 2682 4672 2688 4684
rect 2643 4644 2688 4672
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 4062 4672 4068 4684
rect 4023 4644 4068 4672
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 5810 4672 5816 4684
rect 5771 4644 5816 4672
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 6181 4675 6239 4681
rect 6181 4641 6193 4675
rect 6227 4672 6239 4675
rect 6914 4672 6920 4684
rect 6227 4644 6920 4672
rect 6227 4641 6239 4644
rect 6181 4635 6239 4641
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7300 4681 7328 4712
rect 8386 4700 8392 4712
rect 8444 4700 8450 4752
rect 11701 4743 11759 4749
rect 11701 4709 11713 4743
rect 11747 4740 11759 4743
rect 12434 4740 12440 4752
rect 11747 4712 12440 4740
rect 11747 4709 11759 4712
rect 11701 4703 11759 4709
rect 12434 4700 12440 4712
rect 12492 4700 12498 4752
rect 13541 4743 13599 4749
rect 13541 4740 13553 4743
rect 12544 4712 13553 4740
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4641 7343 4675
rect 8110 4672 8116 4684
rect 8071 4644 8116 4672
rect 7285 4635 7343 4641
rect 8110 4632 8116 4644
rect 8168 4632 8174 4684
rect 8205 4675 8263 4681
rect 8205 4641 8217 4675
rect 8251 4672 8263 4675
rect 12158 4672 12164 4684
rect 8251 4644 12164 4672
rect 8251 4641 8263 4644
rect 8205 4635 8263 4641
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 12544 4672 12572 4712
rect 13541 4709 13553 4712
rect 13587 4709 13599 4743
rect 13541 4703 13599 4709
rect 13630 4700 13636 4752
rect 13688 4740 13694 4752
rect 15304 4749 15332 4780
rect 16206 4768 16212 4820
rect 16264 4808 16270 4820
rect 16942 4808 16948 4820
rect 16264 4780 16948 4808
rect 16264 4768 16270 4780
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 25222 4808 25228 4820
rect 23032 4780 25228 4808
rect 15289 4743 15347 4749
rect 13688 4712 13733 4740
rect 13688 4700 13694 4712
rect 15289 4709 15301 4743
rect 15335 4709 15347 4743
rect 23032 4740 23060 4780
rect 25222 4768 25228 4780
rect 25280 4768 25286 4820
rect 28166 4768 28172 4820
rect 28224 4808 28230 4820
rect 28905 4811 28963 4817
rect 28905 4808 28917 4811
rect 28224 4780 28917 4808
rect 28224 4768 28230 4780
rect 28905 4777 28917 4780
rect 28951 4777 28963 4811
rect 28905 4771 28963 4777
rect 28994 4768 29000 4820
rect 29052 4808 29058 4820
rect 30834 4808 30840 4820
rect 29052 4780 30840 4808
rect 29052 4768 29058 4780
rect 30834 4768 30840 4780
rect 30892 4808 30898 4820
rect 31938 4808 31944 4820
rect 30892 4780 31944 4808
rect 30892 4768 30898 4780
rect 31938 4768 31944 4780
rect 31996 4768 32002 4820
rect 33134 4808 33140 4820
rect 32140 4780 33140 4808
rect 15289 4703 15347 4709
rect 15396 4712 23060 4740
rect 12268 4644 12572 4672
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4573 2651 4607
rect 2593 4567 2651 4573
rect 6273 4607 6331 4613
rect 6273 4573 6285 4607
rect 6319 4604 6331 4607
rect 7098 4604 7104 4616
rect 6319 4576 7104 4604
rect 6319 4573 6331 4576
rect 6273 4567 6331 4573
rect 2608 4536 2636 4567
rect 7098 4564 7104 4576
rect 7156 4564 7162 4616
rect 7374 4604 7380 4616
rect 7335 4576 7380 4604
rect 7374 4564 7380 4576
rect 7432 4564 7438 4616
rect 11609 4607 11667 4613
rect 11609 4573 11621 4607
rect 11655 4604 11667 4607
rect 12069 4607 12127 4613
rect 12069 4604 12081 4607
rect 11655 4576 12081 4604
rect 11655 4573 11667 4576
rect 11609 4567 11667 4573
rect 12069 4573 12081 4576
rect 12115 4604 12127 4607
rect 12268 4604 12296 4644
rect 13170 4632 13176 4684
rect 13228 4672 13234 4684
rect 13449 4675 13507 4681
rect 13449 4672 13461 4675
rect 13228 4644 13461 4672
rect 13228 4632 13234 4644
rect 13449 4641 13461 4644
rect 13495 4641 13507 4675
rect 13449 4635 13507 4641
rect 12115 4576 12296 4604
rect 12115 4573 12127 4576
rect 12069 4567 12127 4573
rect 12802 4564 12808 4616
rect 12860 4604 12866 4616
rect 13265 4607 13323 4613
rect 13265 4604 13277 4607
rect 12860 4576 13277 4604
rect 12860 4564 12866 4576
rect 13265 4573 13277 4576
rect 13311 4573 13323 4607
rect 13265 4567 13323 4573
rect 12434 4536 12440 4548
rect 2608 4508 12440 4536
rect 12434 4496 12440 4508
rect 12492 4496 12498 4548
rect 4154 4468 4160 4480
rect 4115 4440 4160 4468
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 11839 4471 11897 4477
rect 11839 4468 11851 4471
rect 8720 4440 11851 4468
rect 8720 4428 8726 4440
rect 11839 4437 11851 4440
rect 11885 4437 11897 4471
rect 11974 4468 11980 4480
rect 11935 4440 11980 4468
rect 11839 4431 11897 4437
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 13464 4468 13492 4635
rect 13722 4632 13728 4684
rect 13780 4672 13786 4684
rect 15396 4672 15424 4712
rect 23106 4700 23112 4752
rect 23164 4740 23170 4752
rect 24121 4743 24179 4749
rect 24121 4740 24133 4743
rect 23164 4712 24133 4740
rect 23164 4700 23170 4712
rect 24121 4709 24133 4712
rect 24167 4709 24179 4743
rect 25240 4740 25268 4768
rect 26970 4740 26976 4752
rect 25240 4712 26556 4740
rect 24121 4703 24179 4709
rect 13780 4644 15424 4672
rect 13780 4632 13786 4644
rect 16298 4632 16304 4684
rect 16356 4672 16362 4684
rect 17681 4675 17739 4681
rect 17681 4672 17693 4675
rect 16356 4644 17693 4672
rect 16356 4632 16362 4644
rect 17681 4641 17693 4644
rect 17727 4672 17739 4675
rect 18693 4675 18751 4681
rect 18693 4672 18705 4675
rect 17727 4644 18705 4672
rect 17727 4641 17739 4644
rect 17681 4635 17739 4641
rect 18693 4641 18705 4644
rect 18739 4641 18751 4675
rect 18693 4635 18751 4641
rect 19429 4675 19487 4681
rect 19429 4641 19441 4675
rect 19475 4672 19487 4675
rect 20990 4672 20996 4684
rect 19475 4644 20996 4672
rect 19475 4641 19487 4644
rect 19429 4635 19487 4641
rect 20990 4632 20996 4644
rect 21048 4632 21054 4684
rect 22097 4675 22155 4681
rect 22097 4641 22109 4675
rect 22143 4641 22155 4675
rect 22462 4672 22468 4684
rect 22423 4644 22468 4672
rect 22097 4635 22155 4641
rect 13998 4604 14004 4616
rect 13959 4576 14004 4604
rect 13998 4564 14004 4576
rect 14056 4564 14062 4616
rect 15378 4564 15384 4616
rect 15436 4604 15442 4616
rect 15657 4607 15715 4613
rect 15657 4604 15669 4607
rect 15436 4576 15669 4604
rect 15436 4564 15442 4576
rect 15657 4573 15669 4576
rect 15703 4604 15715 4607
rect 16666 4604 16672 4616
rect 15703 4576 16672 4604
rect 15703 4573 15715 4576
rect 15657 4567 15715 4573
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 16850 4604 16856 4616
rect 16811 4576 16856 4604
rect 16850 4564 16856 4576
rect 16908 4564 16914 4616
rect 17405 4607 17463 4613
rect 17405 4573 17417 4607
rect 17451 4573 17463 4607
rect 17862 4604 17868 4616
rect 17823 4576 17868 4604
rect 17405 4567 17463 4573
rect 15746 4536 15752 4548
rect 15442 4508 15752 4536
rect 15442 4477 15470 4508
rect 15746 4496 15752 4508
rect 15804 4496 15810 4548
rect 16022 4496 16028 4548
rect 16080 4536 16086 4548
rect 17420 4536 17448 4567
rect 17862 4564 17868 4576
rect 17920 4564 17926 4616
rect 21910 4604 21916 4616
rect 17972 4576 21916 4604
rect 17972 4536 18000 4576
rect 21910 4564 21916 4576
rect 21968 4564 21974 4616
rect 22112 4604 22140 4635
rect 22462 4632 22468 4644
rect 22520 4632 22526 4684
rect 22738 4672 22744 4684
rect 22699 4644 22744 4672
rect 22738 4632 22744 4644
rect 22796 4632 22802 4684
rect 24581 4675 24639 4681
rect 24581 4641 24593 4675
rect 24627 4641 24639 4675
rect 24854 4672 24860 4684
rect 24815 4644 24860 4672
rect 24581 4635 24639 4641
rect 22554 4604 22560 4616
rect 22112 4576 22560 4604
rect 22554 4564 22560 4576
rect 22612 4604 22618 4616
rect 24302 4604 24308 4616
rect 22612 4576 24308 4604
rect 22612 4564 22618 4576
rect 24302 4564 24308 4576
rect 24360 4564 24366 4616
rect 16080 4508 18000 4536
rect 16080 4496 16086 4508
rect 18230 4496 18236 4548
rect 18288 4536 18294 4548
rect 18785 4539 18843 4545
rect 18785 4536 18797 4539
rect 18288 4508 18797 4536
rect 18288 4496 18294 4508
rect 18785 4505 18797 4508
rect 18831 4505 18843 4539
rect 19242 4536 19248 4548
rect 18785 4499 18843 4505
rect 18892 4508 19248 4536
rect 18892 4480 18920 4508
rect 19242 4496 19248 4508
rect 19300 4496 19306 4548
rect 22189 4539 22247 4545
rect 22189 4505 22201 4539
rect 22235 4536 22247 4539
rect 24026 4536 24032 4548
rect 22235 4508 24032 4536
rect 22235 4505 22247 4508
rect 22189 4499 22247 4505
rect 24026 4496 24032 4508
rect 24084 4536 24090 4548
rect 24596 4536 24624 4635
rect 24854 4632 24860 4644
rect 24912 4632 24918 4684
rect 25041 4675 25099 4681
rect 25041 4641 25053 4675
rect 25087 4641 25099 4675
rect 25041 4635 25099 4641
rect 25225 4675 25283 4681
rect 25225 4641 25237 4675
rect 25271 4672 25283 4675
rect 25406 4672 25412 4684
rect 25271 4644 25412 4672
rect 25271 4641 25283 4644
rect 25225 4635 25283 4641
rect 25056 4604 25084 4635
rect 25406 4632 25412 4644
rect 25464 4632 25470 4684
rect 25501 4675 25559 4681
rect 25501 4641 25513 4675
rect 25547 4672 25559 4675
rect 26418 4672 26424 4684
rect 25547 4644 26424 4672
rect 25547 4641 25559 4644
rect 25501 4635 25559 4641
rect 26418 4632 26424 4644
rect 26476 4632 26482 4684
rect 26528 4681 26556 4712
rect 26620 4712 26976 4740
rect 26620 4681 26648 4712
rect 26970 4700 26976 4712
rect 27028 4700 27034 4752
rect 28261 4743 28319 4749
rect 28261 4709 28273 4743
rect 28307 4740 28319 4743
rect 29086 4740 29092 4752
rect 28307 4712 29092 4740
rect 28307 4709 28319 4712
rect 28261 4703 28319 4709
rect 29086 4700 29092 4712
rect 29144 4700 29150 4752
rect 30193 4743 30251 4749
rect 30193 4709 30205 4743
rect 30239 4740 30251 4743
rect 31110 4740 31116 4752
rect 30239 4712 31116 4740
rect 30239 4709 30251 4712
rect 30193 4703 30251 4709
rect 31110 4700 31116 4712
rect 31168 4700 31174 4752
rect 26513 4675 26571 4681
rect 26513 4641 26525 4675
rect 26559 4641 26571 4675
rect 26513 4635 26571 4641
rect 26605 4675 26663 4681
rect 26605 4641 26617 4675
rect 26651 4641 26663 4675
rect 29178 4672 29184 4684
rect 26605 4635 26663 4641
rect 26712 4644 29184 4672
rect 26712 4604 26740 4644
rect 29178 4632 29184 4644
rect 29236 4672 29242 4684
rect 29730 4672 29736 4684
rect 29236 4644 29736 4672
rect 29236 4632 29242 4644
rect 29730 4632 29736 4644
rect 29788 4632 29794 4684
rect 31018 4672 31024 4684
rect 30979 4644 31024 4672
rect 31018 4632 31024 4644
rect 31076 4632 31082 4684
rect 31205 4675 31263 4681
rect 31205 4641 31217 4675
rect 31251 4672 31263 4675
rect 31938 4672 31944 4684
rect 31251 4644 31944 4672
rect 31251 4641 31263 4644
rect 31205 4635 31263 4641
rect 31938 4632 31944 4644
rect 31996 4632 32002 4684
rect 32030 4632 32036 4684
rect 32088 4672 32094 4684
rect 32140 4681 32168 4780
rect 33134 4768 33140 4780
rect 33192 4808 33198 4820
rect 35069 4811 35127 4817
rect 35069 4808 35081 4811
rect 33192 4780 35081 4808
rect 33192 4768 33198 4780
rect 35069 4777 35081 4780
rect 35115 4777 35127 4811
rect 35069 4771 35127 4777
rect 43625 4811 43683 4817
rect 43625 4777 43637 4811
rect 43671 4808 43683 4811
rect 43714 4808 43720 4820
rect 43671 4780 43720 4808
rect 43671 4777 43683 4780
rect 43625 4771 43683 4777
rect 43714 4768 43720 4780
rect 43772 4768 43778 4820
rect 45557 4811 45615 4817
rect 45557 4777 45569 4811
rect 45603 4808 45615 4811
rect 45738 4808 45744 4820
rect 45603 4780 45744 4808
rect 45603 4777 45615 4780
rect 45557 4771 45615 4777
rect 45738 4768 45744 4780
rect 45796 4768 45802 4820
rect 47872 4780 50384 4808
rect 37182 4740 37188 4752
rect 35176 4712 37188 4740
rect 32125 4675 32183 4681
rect 32125 4672 32137 4675
rect 32088 4644 32137 4672
rect 32088 4632 32094 4644
rect 32125 4641 32137 4644
rect 32171 4641 32183 4675
rect 32125 4635 32183 4641
rect 32401 4675 32459 4681
rect 32401 4641 32413 4675
rect 32447 4672 32459 4675
rect 32490 4672 32496 4684
rect 32447 4644 32496 4672
rect 32447 4641 32459 4644
rect 32401 4635 32459 4641
rect 32490 4632 32496 4644
rect 32548 4632 32554 4684
rect 35176 4681 35204 4712
rect 37182 4700 37188 4712
rect 37240 4700 37246 4752
rect 38102 4700 38108 4752
rect 38160 4740 38166 4752
rect 38160 4712 38516 4740
rect 38160 4700 38166 4712
rect 35161 4675 35219 4681
rect 35161 4641 35173 4675
rect 35207 4641 35219 4675
rect 35161 4635 35219 4641
rect 36265 4675 36323 4681
rect 36265 4641 36277 4675
rect 36311 4641 36323 4675
rect 36265 4635 36323 4641
rect 25056 4576 26740 4604
rect 27065 4607 27123 4613
rect 27065 4573 27077 4607
rect 27111 4573 27123 4607
rect 28626 4604 28632 4616
rect 28587 4576 28632 4604
rect 27065 4567 27123 4573
rect 24084 4508 24624 4536
rect 27080 4536 27108 4567
rect 28626 4564 28632 4576
rect 28684 4564 28690 4616
rect 30558 4564 30564 4616
rect 30616 4604 30622 4616
rect 30745 4607 30803 4613
rect 30745 4604 30757 4607
rect 30616 4576 30757 4604
rect 30616 4564 30622 4576
rect 30745 4573 30757 4576
rect 30791 4573 30803 4607
rect 36078 4604 36084 4616
rect 30745 4567 30803 4573
rect 32140 4576 36084 4604
rect 28537 4539 28595 4545
rect 28537 4536 28549 4539
rect 27080 4508 28549 4536
rect 24084 4496 24090 4508
rect 28537 4505 28549 4508
rect 28583 4505 28595 4539
rect 28537 4499 28595 4505
rect 28902 4496 28908 4548
rect 28960 4536 28966 4548
rect 32140 4536 32168 4576
rect 36078 4564 36084 4576
rect 36136 4604 36142 4616
rect 36280 4604 36308 4635
rect 36354 4632 36360 4684
rect 36412 4672 36418 4684
rect 36449 4675 36507 4681
rect 36449 4672 36461 4675
rect 36412 4644 36461 4672
rect 36412 4632 36418 4644
rect 36449 4641 36461 4644
rect 36495 4641 36507 4675
rect 38378 4672 38384 4684
rect 38339 4644 38384 4672
rect 36449 4635 36507 4641
rect 38378 4632 38384 4644
rect 38436 4632 38442 4684
rect 38488 4681 38516 4712
rect 40034 4700 40040 4752
rect 40092 4740 40098 4752
rect 40092 4712 43576 4740
rect 40092 4700 40098 4712
rect 38473 4675 38531 4681
rect 38473 4641 38485 4675
rect 38519 4641 38531 4675
rect 38473 4635 38531 4641
rect 38930 4632 38936 4684
rect 38988 4672 38994 4684
rect 41141 4675 41199 4681
rect 41141 4672 41153 4675
rect 38988 4644 41153 4672
rect 38988 4632 38994 4644
rect 41141 4641 41153 4644
rect 41187 4641 41199 4675
rect 41141 4635 41199 4641
rect 41371 4675 41429 4681
rect 41371 4641 41383 4675
rect 41417 4672 41429 4675
rect 41966 4672 41972 4684
rect 41417 4644 41972 4672
rect 41417 4641 41429 4644
rect 41371 4635 41429 4641
rect 41966 4632 41972 4644
rect 42024 4632 42030 4684
rect 43548 4681 43576 4712
rect 43349 4675 43407 4681
rect 43349 4672 43361 4675
rect 42076 4644 43361 4672
rect 36136 4576 36308 4604
rect 36136 4564 36142 4576
rect 35342 4536 35348 4548
rect 28960 4508 32168 4536
rect 35303 4508 35348 4536
rect 28960 4496 28966 4508
rect 35342 4496 35348 4508
rect 35400 4496 35406 4548
rect 36280 4536 36308 4576
rect 36817 4607 36875 4613
rect 36817 4573 36829 4607
rect 36863 4604 36875 4607
rect 37274 4604 37280 4616
rect 36863 4576 37280 4604
rect 36863 4573 36875 4576
rect 36817 4567 36875 4573
rect 37274 4564 37280 4576
rect 37332 4564 37338 4616
rect 40589 4607 40647 4613
rect 40589 4573 40601 4607
rect 40635 4604 40647 4607
rect 40862 4604 40868 4616
rect 40635 4576 40868 4604
rect 40635 4573 40647 4576
rect 40589 4567 40647 4573
rect 40862 4564 40868 4576
rect 40920 4564 40926 4616
rect 41230 4564 41236 4616
rect 41288 4604 41294 4616
rect 41601 4607 41659 4613
rect 41601 4604 41613 4607
rect 41288 4576 41613 4604
rect 41288 4564 41294 4576
rect 41601 4573 41613 4576
rect 41647 4573 41659 4607
rect 41601 4567 41659 4573
rect 37826 4536 37832 4548
rect 36280 4508 37832 4536
rect 37826 4496 37832 4508
rect 37884 4496 37890 4548
rect 40402 4496 40408 4548
rect 40460 4536 40466 4548
rect 42076 4536 42104 4644
rect 43349 4641 43361 4644
rect 43395 4641 43407 4675
rect 43349 4635 43407 4641
rect 43533 4675 43591 4681
rect 43533 4641 43545 4675
rect 43579 4641 43591 4675
rect 43533 4635 43591 4641
rect 45373 4675 45431 4681
rect 45373 4641 45385 4675
rect 45419 4672 45431 4675
rect 45462 4672 45468 4684
rect 45419 4644 45468 4672
rect 45419 4641 45431 4644
rect 45373 4635 45431 4641
rect 43548 4604 43576 4635
rect 45462 4632 45468 4644
rect 45520 4632 45526 4684
rect 46566 4672 46572 4684
rect 46527 4644 46572 4672
rect 46566 4632 46572 4644
rect 46624 4632 46630 4684
rect 47872 4681 47900 4780
rect 47946 4700 47952 4752
rect 48004 4740 48010 4752
rect 50356 4740 50384 4780
rect 50430 4768 50436 4820
rect 50488 4808 50494 4820
rect 50488 4780 52132 4808
rect 50488 4768 50494 4780
rect 50617 4743 50675 4749
rect 50617 4740 50629 4743
rect 48004 4712 48049 4740
rect 50356 4712 50629 4740
rect 48004 4700 48010 4712
rect 50617 4709 50629 4712
rect 50663 4740 50675 4743
rect 50798 4740 50804 4752
rect 50663 4712 50804 4740
rect 50663 4709 50675 4712
rect 50617 4703 50675 4709
rect 50798 4700 50804 4712
rect 50856 4700 50862 4752
rect 47857 4675 47915 4681
rect 47857 4641 47869 4675
rect 47903 4641 47915 4675
rect 47857 4635 47915 4641
rect 48961 4675 49019 4681
rect 48961 4641 48973 4675
rect 49007 4672 49019 4675
rect 49050 4672 49056 4684
rect 49007 4644 49056 4672
rect 49007 4641 49019 4644
rect 48961 4635 49019 4641
rect 49050 4632 49056 4644
rect 49108 4672 49114 4684
rect 51718 4672 51724 4684
rect 49108 4644 51724 4672
rect 49108 4632 49114 4644
rect 51718 4632 51724 4644
rect 51776 4632 51782 4684
rect 52104 4681 52132 4780
rect 58618 4768 58624 4820
rect 58676 4808 58682 4820
rect 58802 4808 58808 4820
rect 58676 4780 58808 4808
rect 58676 4768 58682 4780
rect 58802 4768 58808 4780
rect 58860 4768 58866 4820
rect 55769 4743 55827 4749
rect 55769 4709 55781 4743
rect 55815 4740 55827 4743
rect 57606 4740 57612 4752
rect 55815 4712 57612 4740
rect 55815 4709 55827 4712
rect 55769 4703 55827 4709
rect 57606 4700 57612 4712
rect 57664 4700 57670 4752
rect 60182 4740 60188 4752
rect 58636 4712 60188 4740
rect 52089 4675 52147 4681
rect 52089 4641 52101 4675
rect 52135 4641 52147 4675
rect 52454 4672 52460 4684
rect 52415 4644 52460 4672
rect 52089 4635 52147 4641
rect 52454 4632 52460 4644
rect 52512 4632 52518 4684
rect 56318 4632 56324 4684
rect 56376 4681 56382 4684
rect 56376 4675 56425 4681
rect 56376 4641 56379 4675
rect 56413 4641 56425 4675
rect 56502 4672 56508 4684
rect 56463 4644 56508 4672
rect 56376 4635 56425 4641
rect 56376 4632 56382 4635
rect 56502 4632 56508 4644
rect 56560 4672 56566 4684
rect 58636 4672 58664 4712
rect 60182 4700 60188 4712
rect 60240 4700 60246 4752
rect 58802 4672 58808 4684
rect 56560 4644 58664 4672
rect 58763 4644 58808 4672
rect 56560 4632 56566 4644
rect 58802 4632 58808 4644
rect 58860 4632 58866 4684
rect 46477 4607 46535 4613
rect 46477 4604 46489 4607
rect 43548 4576 46489 4604
rect 46477 4573 46489 4576
rect 46523 4573 46535 4607
rect 46477 4567 46535 4573
rect 47029 4607 47087 4613
rect 47029 4573 47041 4607
rect 47075 4604 47087 4607
rect 48774 4604 48780 4616
rect 47075 4576 48780 4604
rect 47075 4573 47087 4576
rect 47029 4567 47087 4573
rect 48774 4564 48780 4576
rect 48832 4564 48838 4616
rect 49237 4607 49295 4613
rect 49237 4573 49249 4607
rect 49283 4604 49295 4607
rect 49418 4604 49424 4616
rect 49283 4576 49424 4604
rect 49283 4573 49295 4576
rect 49237 4567 49295 4573
rect 49418 4564 49424 4576
rect 49476 4564 49482 4616
rect 50430 4564 50436 4616
rect 50488 4604 50494 4616
rect 51445 4607 51503 4613
rect 51445 4604 51457 4607
rect 50488 4576 51457 4604
rect 50488 4564 50494 4576
rect 51445 4573 51457 4576
rect 51491 4573 51503 4607
rect 51445 4567 51503 4573
rect 52181 4607 52239 4613
rect 52181 4573 52193 4607
rect 52227 4573 52239 4607
rect 52181 4567 52239 4573
rect 40460 4508 42104 4536
rect 52196 4536 52224 4567
rect 52270 4564 52276 4616
rect 52328 4604 52334 4616
rect 52365 4607 52423 4613
rect 52365 4604 52377 4607
rect 52328 4576 52377 4604
rect 52328 4564 52334 4576
rect 52365 4573 52377 4576
rect 52411 4573 52423 4607
rect 52365 4567 52423 4573
rect 55677 4607 55735 4613
rect 55677 4573 55689 4607
rect 55723 4573 55735 4607
rect 57974 4604 57980 4616
rect 57935 4576 57980 4604
rect 55677 4567 55735 4573
rect 55398 4536 55404 4548
rect 52196 4508 55404 4536
rect 40460 4496 40466 4508
rect 55398 4496 55404 4508
rect 55456 4536 55462 4548
rect 55692 4536 55720 4567
rect 57974 4564 57980 4576
rect 58032 4564 58038 4616
rect 58989 4607 59047 4613
rect 58989 4604 59001 4607
rect 58084 4576 59001 4604
rect 55456 4508 55720 4536
rect 55456 4496 55462 4508
rect 56686 4496 56692 4548
rect 56744 4536 56750 4548
rect 58084 4536 58112 4576
rect 58989 4573 59001 4576
rect 59035 4573 59047 4607
rect 58989 4567 59047 4573
rect 58434 4536 58440 4548
rect 56744 4508 58112 4536
rect 58395 4508 58440 4536
rect 56744 4496 56750 4508
rect 58434 4496 58440 4508
rect 58492 4496 58498 4548
rect 15427 4471 15485 4477
rect 15427 4468 15439 4471
rect 13464 4440 15439 4468
rect 15427 4437 15439 4440
rect 15473 4437 15485 4471
rect 15427 4431 15485 4437
rect 15562 4428 15568 4480
rect 15620 4468 15626 4480
rect 15933 4471 15991 4477
rect 15620 4440 15665 4468
rect 15620 4428 15626 4440
rect 15933 4437 15945 4471
rect 15979 4468 15991 4471
rect 18874 4468 18880 4480
rect 15979 4440 18880 4468
rect 15979 4437 15991 4440
rect 15933 4431 15991 4437
rect 18874 4428 18880 4440
rect 18932 4428 18938 4480
rect 18966 4428 18972 4480
rect 19024 4468 19030 4480
rect 20346 4468 20352 4480
rect 19024 4440 20352 4468
rect 19024 4428 19030 4440
rect 20346 4428 20352 4440
rect 20404 4428 20410 4480
rect 28350 4428 28356 4480
rect 28408 4477 28414 4480
rect 28408 4471 28457 4477
rect 28408 4437 28411 4471
rect 28445 4437 28457 4471
rect 28408 4431 28457 4437
rect 28408 4428 28414 4431
rect 28718 4428 28724 4480
rect 28776 4468 28782 4480
rect 31018 4468 31024 4480
rect 28776 4440 31024 4468
rect 28776 4428 28782 4440
rect 31018 4428 31024 4440
rect 31076 4428 31082 4480
rect 31294 4428 31300 4480
rect 31352 4468 31358 4480
rect 32030 4468 32036 4480
rect 31352 4440 32036 4468
rect 31352 4428 31358 4440
rect 32030 4428 32036 4440
rect 32088 4428 32094 4480
rect 33318 4428 33324 4480
rect 33376 4468 33382 4480
rect 33689 4471 33747 4477
rect 33689 4468 33701 4471
rect 33376 4440 33701 4468
rect 33376 4428 33382 4440
rect 33689 4437 33701 4440
rect 33735 4468 33747 4471
rect 34974 4468 34980 4480
rect 33735 4440 34980 4468
rect 33735 4437 33747 4440
rect 33689 4431 33747 4437
rect 34974 4428 34980 4440
rect 35032 4428 35038 4480
rect 35069 4471 35127 4477
rect 35069 4437 35081 4471
rect 35115 4468 35127 4471
rect 37458 4468 37464 4480
rect 35115 4440 37464 4468
rect 35115 4437 35127 4440
rect 35069 4431 35127 4437
rect 37458 4428 37464 4440
rect 37516 4428 37522 4480
rect 38102 4428 38108 4480
rect 38160 4468 38166 4480
rect 38197 4471 38255 4477
rect 38197 4468 38209 4471
rect 38160 4440 38209 4468
rect 38160 4428 38166 4440
rect 38197 4437 38209 4440
rect 38243 4437 38255 4471
rect 38654 4468 38660 4480
rect 38615 4440 38660 4468
rect 38197 4431 38255 4437
rect 38654 4428 38660 4440
rect 38712 4428 38718 4480
rect 46934 4428 46940 4480
rect 46992 4468 46998 4480
rect 55674 4468 55680 4480
rect 46992 4440 55680 4468
rect 46992 4428 46998 4440
rect 55674 4428 55680 4440
rect 55732 4428 55738 4480
rect 1104 4378 62192 4400
rect 1104 4326 11163 4378
rect 11215 4326 11227 4378
rect 11279 4326 11291 4378
rect 11343 4326 11355 4378
rect 11407 4326 31526 4378
rect 31578 4326 31590 4378
rect 31642 4326 31654 4378
rect 31706 4326 31718 4378
rect 31770 4326 51888 4378
rect 51940 4326 51952 4378
rect 52004 4326 52016 4378
rect 52068 4326 52080 4378
rect 52132 4326 62192 4378
rect 1104 4304 62192 4326
rect 6914 4224 6920 4276
rect 6972 4264 6978 4276
rect 8018 4264 8024 4276
rect 6972 4236 8024 4264
rect 6972 4224 6978 4236
rect 8018 4224 8024 4236
rect 8076 4264 8082 4276
rect 11974 4264 11980 4276
rect 8076 4236 11980 4264
rect 8076 4224 8082 4236
rect 11974 4224 11980 4236
rect 12032 4264 12038 4276
rect 13630 4264 13636 4276
rect 12032 4236 13636 4264
rect 12032 4224 12038 4236
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 22462 4264 22468 4276
rect 14056 4236 22468 4264
rect 14056 4224 14062 4236
rect 22462 4224 22468 4236
rect 22520 4224 22526 4276
rect 27798 4224 27804 4276
rect 27856 4264 27862 4276
rect 28902 4264 28908 4276
rect 27856 4236 28908 4264
rect 27856 4224 27862 4236
rect 28902 4224 28908 4236
rect 28960 4224 28966 4276
rect 29917 4267 29975 4273
rect 29917 4233 29929 4267
rect 29963 4264 29975 4267
rect 31386 4264 31392 4276
rect 29963 4236 31392 4264
rect 29963 4233 29975 4236
rect 29917 4227 29975 4233
rect 31386 4224 31392 4236
rect 31444 4264 31450 4276
rect 32214 4264 32220 4276
rect 31444 4236 32220 4264
rect 31444 4224 31450 4236
rect 32214 4224 32220 4236
rect 32272 4224 32278 4276
rect 33042 4224 33048 4276
rect 33100 4264 33106 4276
rect 35069 4267 35127 4273
rect 35069 4264 35081 4267
rect 33100 4236 35081 4264
rect 33100 4224 33106 4236
rect 35069 4233 35081 4236
rect 35115 4264 35127 4267
rect 37366 4264 37372 4276
rect 35115 4236 37372 4264
rect 35115 4233 35127 4236
rect 35069 4227 35127 4233
rect 37366 4224 37372 4236
rect 37424 4224 37430 4276
rect 41046 4224 41052 4276
rect 41104 4264 41110 4276
rect 43993 4267 44051 4273
rect 43993 4264 44005 4267
rect 41104 4236 44005 4264
rect 41104 4224 41110 4236
rect 43993 4233 44005 4236
rect 44039 4264 44051 4267
rect 46842 4264 46848 4276
rect 44039 4236 46848 4264
rect 44039 4233 44051 4236
rect 43993 4227 44051 4233
rect 46842 4224 46848 4236
rect 46900 4224 46906 4276
rect 49694 4224 49700 4276
rect 49752 4264 49758 4276
rect 51350 4264 51356 4276
rect 49752 4236 51356 4264
rect 49752 4224 49758 4236
rect 51350 4224 51356 4236
rect 51408 4264 51414 4276
rect 52270 4264 52276 4276
rect 51408 4236 52276 4264
rect 51408 4224 51414 4236
rect 52270 4224 52276 4236
rect 52328 4224 52334 4276
rect 6822 4156 6828 4208
rect 6880 4196 6886 4208
rect 6880 4168 9168 4196
rect 6880 4156 6886 4168
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4128 3203 4131
rect 4522 4128 4528 4140
rect 3191 4100 4384 4128
rect 4483 4100 4528 4128
rect 3191 4097 3203 4100
rect 3145 4091 3203 4097
rect 2593 4063 2651 4069
rect 2593 4029 2605 4063
rect 2639 4029 2651 4063
rect 2593 4023 2651 4029
rect 2608 3924 2636 4023
rect 2682 4020 2688 4072
rect 2740 4060 2746 4072
rect 3970 4060 3976 4072
rect 2740 4032 2833 4060
rect 3931 4032 3976 4060
rect 2740 4020 2746 4032
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 4065 4063 4123 4069
rect 4065 4029 4077 4063
rect 4111 4029 4123 4063
rect 4356 4060 4384 4100
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 7190 4128 7196 4140
rect 5184 4100 7196 4128
rect 5184 4060 5212 4100
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 7742 4128 7748 4140
rect 7703 4100 7748 4128
rect 7742 4088 7748 4100
rect 7800 4128 7806 4140
rect 9030 4128 9036 4140
rect 7800 4100 9036 4128
rect 7800 4088 7806 4100
rect 9030 4088 9036 4100
rect 9088 4088 9094 4140
rect 9140 4128 9168 4168
rect 11054 4156 11060 4208
rect 11112 4196 11118 4208
rect 11606 4196 11612 4208
rect 11112 4168 11612 4196
rect 11112 4156 11118 4168
rect 11606 4156 11612 4168
rect 11664 4196 11670 4208
rect 19978 4196 19984 4208
rect 11664 4168 19984 4196
rect 11664 4156 11670 4168
rect 19978 4156 19984 4168
rect 20036 4156 20042 4208
rect 25884 4168 28396 4196
rect 13538 4128 13544 4140
rect 9140 4100 13544 4128
rect 13188 4072 13216 4100
rect 13538 4088 13544 4100
rect 13596 4088 13602 4140
rect 15194 4128 15200 4140
rect 14108 4100 15200 4128
rect 5350 4060 5356 4072
rect 4356 4032 5212 4060
rect 5311 4032 5356 4060
rect 4065 4023 4123 4029
rect 2700 3992 2728 4020
rect 4080 3992 4108 4023
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 5445 4063 5503 4069
rect 5445 4029 5457 4063
rect 5491 4060 5503 4063
rect 5718 4060 5724 4072
rect 5491 4032 5724 4060
rect 5491 4029 5503 4032
rect 5445 4023 5503 4029
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 5905 4063 5963 4069
rect 5905 4029 5917 4063
rect 5951 4060 5963 4063
rect 7285 4063 7343 4069
rect 7285 4060 7297 4063
rect 5951 4032 7297 4060
rect 5951 4029 5963 4032
rect 5905 4023 5963 4029
rect 7285 4029 7297 4032
rect 7331 4029 7343 4063
rect 7466 4060 7472 4072
rect 7427 4032 7472 4060
rect 7285 4023 7343 4029
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 7837 4063 7895 4069
rect 7837 4029 7849 4063
rect 7883 4029 7895 4063
rect 7837 4023 7895 4029
rect 8849 4063 8907 4069
rect 8849 4029 8861 4063
rect 8895 4029 8907 4063
rect 8849 4023 8907 4029
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4029 13139 4063
rect 13081 4023 13139 4029
rect 7558 3992 7564 4004
rect 2700 3964 7564 3992
rect 7558 3952 7564 3964
rect 7616 3952 7622 4004
rect 6730 3924 6736 3936
rect 2608 3896 6736 3924
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 6914 3924 6920 3936
rect 6875 3896 6920 3924
rect 6914 3884 6920 3896
rect 6972 3884 6978 3936
rect 7852 3924 7880 4023
rect 8662 3952 8668 4004
rect 8720 3992 8726 4004
rect 8864 3992 8892 4023
rect 9950 3992 9956 4004
rect 8720 3964 8892 3992
rect 8956 3964 9956 3992
rect 8720 3952 8726 3964
rect 8956 3924 8984 3964
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 13096 3992 13124 4023
rect 13170 4020 13176 4072
rect 13228 4060 13234 4072
rect 14108 4060 14136 4100
rect 15194 4088 15200 4100
rect 15252 4088 15258 4140
rect 18230 4128 18236 4140
rect 18191 4100 18236 4128
rect 18230 4088 18236 4100
rect 18288 4088 18294 4140
rect 20162 4128 20168 4140
rect 20123 4100 20168 4128
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 22554 4088 22560 4140
rect 22612 4128 22618 4140
rect 24854 4128 24860 4140
rect 22612 4100 24860 4128
rect 22612 4088 22618 4100
rect 24854 4088 24860 4100
rect 24912 4088 24918 4140
rect 25685 4131 25743 4137
rect 25685 4097 25697 4131
rect 25731 4128 25743 4131
rect 25884 4128 25912 4168
rect 28258 4128 28264 4140
rect 25731 4100 25912 4128
rect 25976 4100 28264 4128
rect 25731 4097 25743 4100
rect 25685 4091 25743 4097
rect 13228 4032 13273 4060
rect 13372 4032 14136 4060
rect 13228 4020 13234 4032
rect 13262 3992 13268 4004
rect 13096 3964 13268 3992
rect 13262 3952 13268 3964
rect 13320 3992 13326 4004
rect 13372 3992 13400 4032
rect 14182 4020 14188 4072
rect 14240 4060 14246 4072
rect 14921 4063 14979 4069
rect 14921 4060 14933 4063
rect 14240 4032 14933 4060
rect 14240 4020 14246 4032
rect 14921 4029 14933 4032
rect 14967 4029 14979 4063
rect 15286 4060 15292 4072
rect 15247 4032 15292 4060
rect 14921 4023 14979 4029
rect 15286 4020 15292 4032
rect 15344 4020 15350 4072
rect 16666 4060 16672 4072
rect 16627 4032 16672 4060
rect 16666 4020 16672 4032
rect 16724 4020 16730 4072
rect 16850 4020 16856 4072
rect 16908 4060 16914 4072
rect 16945 4063 17003 4069
rect 16945 4060 16957 4063
rect 16908 4032 16957 4060
rect 16908 4020 16914 4032
rect 16945 4029 16957 4032
rect 16991 4029 17003 4063
rect 16945 4023 17003 4029
rect 17129 4063 17187 4069
rect 17129 4029 17141 4063
rect 17175 4060 17187 4063
rect 17218 4060 17224 4072
rect 17175 4032 17224 4060
rect 17175 4029 17187 4032
rect 17129 4023 17187 4029
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 18782 4020 18788 4072
rect 18840 4060 18846 4072
rect 19058 4069 19064 4072
rect 18923 4063 18981 4069
rect 18923 4060 18935 4063
rect 18840 4032 18935 4060
rect 18840 4020 18846 4032
rect 18923 4029 18935 4032
rect 18969 4029 18981 4063
rect 18923 4023 18981 4029
rect 19049 4063 19064 4069
rect 19049 4029 19061 4063
rect 19049 4023 19064 4029
rect 19058 4020 19064 4023
rect 19116 4020 19122 4072
rect 19242 4020 19248 4072
rect 19300 4020 19306 4072
rect 20070 4060 20076 4072
rect 20031 4032 20076 4060
rect 20070 4020 20076 4032
rect 20128 4020 20134 4072
rect 20346 4060 20352 4072
rect 20307 4032 20352 4060
rect 20346 4020 20352 4032
rect 20404 4020 20410 4072
rect 22465 4063 22523 4069
rect 22465 4029 22477 4063
rect 22511 4060 22523 4063
rect 22511 4032 23336 4060
rect 22511 4029 22523 4032
rect 22465 4023 22523 4029
rect 13320 3964 13400 3992
rect 13320 3952 13326 3964
rect 13446 3952 13452 4004
rect 13504 3992 13510 4004
rect 13633 3995 13691 4001
rect 13633 3992 13645 3995
rect 13504 3964 13645 3992
rect 13504 3952 13510 3964
rect 13633 3961 13645 3964
rect 13679 3961 13691 3995
rect 13633 3955 13691 3961
rect 14737 3995 14795 4001
rect 14737 3961 14749 3995
rect 14783 3992 14795 3995
rect 16022 3992 16028 4004
rect 14783 3964 16028 3992
rect 14783 3961 14795 3964
rect 14737 3955 14795 3961
rect 16022 3952 16028 3964
rect 16080 3952 16086 4004
rect 16117 3995 16175 4001
rect 16117 3961 16129 3995
rect 16163 3961 16175 3995
rect 18322 3992 18328 4004
rect 18283 3964 18328 3992
rect 16117 3955 16175 3961
rect 7852 3896 8984 3924
rect 9033 3927 9091 3933
rect 9033 3893 9045 3927
rect 9079 3924 9091 3927
rect 9122 3924 9128 3936
rect 9079 3896 9128 3924
rect 9079 3893 9091 3896
rect 9033 3887 9091 3893
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 16132 3924 16160 3955
rect 18322 3952 18328 3964
rect 18380 3952 18386 4004
rect 19260 3992 19288 4020
rect 23308 4004 23336 4032
rect 23658 4020 23664 4072
rect 23716 4060 23722 4072
rect 23753 4063 23811 4069
rect 23753 4060 23765 4063
rect 23716 4032 23765 4060
rect 23716 4020 23722 4032
rect 23753 4029 23765 4032
rect 23799 4029 23811 4063
rect 23753 4023 23811 4029
rect 23842 4020 23848 4072
rect 23900 4060 23906 4072
rect 25976 4069 26004 4100
rect 28258 4088 28264 4100
rect 28316 4088 28322 4140
rect 28368 4128 28396 4168
rect 34974 4156 34980 4208
rect 35032 4196 35038 4208
rect 37734 4196 37740 4208
rect 35032 4168 37740 4196
rect 35032 4156 35038 4168
rect 37734 4156 37740 4168
rect 37792 4156 37798 4208
rect 38856 4168 40172 4196
rect 31202 4128 31208 4140
rect 28368 4100 31208 4128
rect 31202 4088 31208 4100
rect 31260 4128 31266 4140
rect 37001 4131 37059 4137
rect 37001 4128 37013 4131
rect 31260 4100 37013 4128
rect 31260 4088 31266 4100
rect 37001 4097 37013 4100
rect 37047 4097 37059 4131
rect 37001 4091 37059 4097
rect 37108 4100 37412 4128
rect 25961 4063 26019 4069
rect 23900 4032 23945 4060
rect 23900 4020 23906 4032
rect 25961 4029 25973 4063
rect 26007 4029 26019 4063
rect 25961 4023 26019 4029
rect 26050 4020 26056 4072
rect 26108 4060 26114 4072
rect 26145 4063 26203 4069
rect 26145 4060 26157 4063
rect 26108 4032 26157 4060
rect 26108 4020 26114 4032
rect 26145 4029 26157 4032
rect 26191 4060 26203 4063
rect 27157 4063 27215 4069
rect 27157 4060 27169 4063
rect 26191 4032 27169 4060
rect 26191 4029 26203 4032
rect 26145 4023 26203 4029
rect 27157 4029 27169 4032
rect 27203 4029 27215 4063
rect 28994 4060 29000 4072
rect 27157 4023 27215 4029
rect 27264 4032 29000 4060
rect 20806 3992 20812 4004
rect 19260 3964 20812 3992
rect 20806 3952 20812 3964
rect 20864 3952 20870 4004
rect 23290 3952 23296 4004
rect 23348 3992 23354 4004
rect 24305 3995 24363 4001
rect 24305 3992 24317 3995
rect 23348 3964 24317 3992
rect 23348 3952 23354 3964
rect 24305 3961 24317 3964
rect 24351 3961 24363 3995
rect 24305 3955 24363 3961
rect 25133 3995 25191 4001
rect 25133 3961 25145 3995
rect 25179 3992 25191 3995
rect 26786 3992 26792 4004
rect 25179 3964 26792 3992
rect 25179 3961 25191 3964
rect 25133 3955 25191 3961
rect 26786 3952 26792 3964
rect 26844 3952 26850 4004
rect 26973 3995 27031 4001
rect 26973 3961 26985 3995
rect 27019 3992 27031 3995
rect 27264 3992 27292 4032
rect 28994 4020 29000 4032
rect 29052 4020 29058 4072
rect 29270 4020 29276 4072
rect 29328 4060 29334 4072
rect 29546 4060 29552 4072
rect 29328 4032 29552 4060
rect 29328 4020 29334 4032
rect 29546 4020 29552 4032
rect 29604 4020 29610 4072
rect 30193 4063 30251 4069
rect 30193 4029 30205 4063
rect 30239 4060 30251 4063
rect 31018 4060 31024 4072
rect 30239 4032 31024 4060
rect 30239 4029 30251 4032
rect 30193 4023 30251 4029
rect 31018 4020 31024 4032
rect 31076 4020 31082 4072
rect 31294 4020 31300 4072
rect 31352 4060 31358 4072
rect 31481 4063 31539 4069
rect 31481 4060 31493 4063
rect 31352 4032 31493 4060
rect 31352 4020 31358 4032
rect 31481 4029 31493 4032
rect 31527 4029 31539 4063
rect 31757 4063 31815 4069
rect 31757 4060 31769 4063
rect 31481 4023 31539 4029
rect 31588 4032 31769 4060
rect 30098 3992 30104 4004
rect 27019 3964 27292 3992
rect 30059 3964 30104 3992
rect 27019 3961 27031 3964
rect 26973 3955 27031 3961
rect 30098 3952 30104 3964
rect 30156 3952 30162 4004
rect 30653 3995 30711 4001
rect 30653 3961 30665 3995
rect 30699 3992 30711 3995
rect 30926 3992 30932 4004
rect 30699 3964 30932 3992
rect 30699 3961 30711 3964
rect 30653 3955 30711 3961
rect 30926 3952 30932 3964
rect 30984 3952 30990 4004
rect 31110 3952 31116 4004
rect 31168 3992 31174 4004
rect 31588 3992 31616 4032
rect 31757 4029 31769 4032
rect 31803 4029 31815 4063
rect 31757 4023 31815 4029
rect 34885 4063 34943 4069
rect 34885 4029 34897 4063
rect 34931 4060 34943 4063
rect 34974 4060 34980 4072
rect 34931 4032 34980 4060
rect 34931 4029 34943 4032
rect 34885 4023 34943 4029
rect 34974 4020 34980 4032
rect 35032 4020 35038 4072
rect 35989 4063 36047 4069
rect 35989 4029 36001 4063
rect 36035 4060 36047 4063
rect 36078 4060 36084 4072
rect 36035 4032 36084 4060
rect 36035 4029 36047 4032
rect 35989 4023 36047 4029
rect 36078 4020 36084 4032
rect 36136 4020 36142 4072
rect 37108 4060 37136 4100
rect 37274 4060 37280 4072
rect 36188 4032 37136 4060
rect 37235 4032 37280 4060
rect 31168 3964 31616 3992
rect 31168 3952 31174 3964
rect 32490 3952 32496 4004
rect 32548 3992 32554 4004
rect 36188 3992 36216 4032
rect 37274 4020 37280 4032
rect 37332 4020 37338 4072
rect 37384 4060 37412 4100
rect 37458 4088 37464 4140
rect 37516 4128 37522 4140
rect 37918 4128 37924 4140
rect 37516 4100 37924 4128
rect 37516 4088 37522 4100
rect 37918 4088 37924 4100
rect 37976 4128 37982 4140
rect 38562 4128 38568 4140
rect 37976 4100 38568 4128
rect 37976 4088 37982 4100
rect 38562 4088 38568 4100
rect 38620 4128 38626 4140
rect 38856 4128 38884 4168
rect 38620 4100 38884 4128
rect 38620 4088 38626 4100
rect 38930 4088 38936 4140
rect 38988 4128 38994 4140
rect 39117 4131 39175 4137
rect 39117 4128 39129 4131
rect 38988 4100 39129 4128
rect 38988 4088 38994 4100
rect 39117 4097 39129 4100
rect 39163 4097 39175 4131
rect 40034 4128 40040 4140
rect 39117 4091 39175 4097
rect 39224 4100 40040 4128
rect 39224 4060 39252 4100
rect 40034 4088 40040 4100
rect 40092 4088 40098 4140
rect 40144 4128 40172 4168
rect 45738 4156 45744 4208
rect 45796 4196 45802 4208
rect 49418 4196 49424 4208
rect 45796 4168 49280 4196
rect 49379 4168 49424 4196
rect 45796 4156 45802 4168
rect 40494 4128 40500 4140
rect 40144 4100 40500 4128
rect 40494 4088 40500 4100
rect 40552 4128 40558 4140
rect 40589 4131 40647 4137
rect 40589 4128 40601 4131
rect 40552 4100 40601 4128
rect 40552 4088 40558 4100
rect 40589 4097 40601 4100
rect 40635 4097 40647 4131
rect 40862 4128 40868 4140
rect 40823 4100 40868 4128
rect 40589 4091 40647 4097
rect 40862 4088 40868 4100
rect 40920 4088 40926 4140
rect 45554 4088 45560 4140
rect 45612 4128 45618 4140
rect 47029 4131 47087 4137
rect 47029 4128 47041 4131
rect 45612 4100 47041 4128
rect 45612 4088 45618 4100
rect 47029 4097 47041 4100
rect 47075 4097 47087 4131
rect 49252 4128 49280 4168
rect 49418 4156 49424 4168
rect 49476 4156 49482 4208
rect 49252 4100 49648 4128
rect 47029 4091 47087 4097
rect 37384 4032 39252 4060
rect 39298 4020 39304 4072
rect 39356 4060 39362 4072
rect 39393 4063 39451 4069
rect 39393 4060 39405 4063
rect 39356 4032 39405 4060
rect 39356 4020 39362 4032
rect 39393 4029 39405 4032
rect 39439 4029 39451 4063
rect 39574 4060 39580 4072
rect 39535 4032 39580 4060
rect 39393 4023 39451 4029
rect 39574 4020 39580 4032
rect 39632 4020 39638 4072
rect 43070 4020 43076 4072
rect 43128 4060 43134 4072
rect 43809 4063 43867 4069
rect 43809 4060 43821 4063
rect 43128 4032 43821 4060
rect 43128 4020 43134 4032
rect 43809 4029 43821 4032
rect 43855 4029 43867 4063
rect 44910 4060 44916 4072
rect 44871 4032 44916 4060
rect 43809 4023 43867 4029
rect 32548 3964 36216 3992
rect 32548 3952 32554 3964
rect 36630 3952 36636 4004
rect 36688 3992 36694 4004
rect 37185 3995 37243 4001
rect 37185 3992 37197 3995
rect 36688 3964 37197 3992
rect 36688 3952 36694 3964
rect 37185 3961 37197 3964
rect 37231 3961 37243 3995
rect 37185 3955 37243 3961
rect 37737 3995 37795 4001
rect 37737 3961 37749 3995
rect 37783 3992 37795 3995
rect 38194 3992 38200 4004
rect 37783 3964 38200 3992
rect 37783 3961 37795 3964
rect 37737 3955 37795 3961
rect 38194 3952 38200 3964
rect 38252 3952 38258 4004
rect 38565 3995 38623 4001
rect 38565 3961 38577 3995
rect 38611 3992 38623 3995
rect 39206 3992 39212 4004
rect 38611 3964 39212 3992
rect 38611 3961 38623 3964
rect 38565 3955 38623 3961
rect 39206 3952 39212 3964
rect 39264 3952 39270 4004
rect 43824 3992 43852 4023
rect 44910 4020 44916 4032
rect 44968 4020 44974 4072
rect 45462 4020 45468 4072
rect 45520 4060 45526 4072
rect 47121 4063 47179 4069
rect 47121 4060 47133 4063
rect 45520 4032 47133 4060
rect 45520 4020 45526 4032
rect 47121 4029 47133 4032
rect 47167 4029 47179 4063
rect 47121 4023 47179 4029
rect 47489 4063 47547 4069
rect 47489 4029 47501 4063
rect 47535 4060 47547 4063
rect 47578 4060 47584 4072
rect 47535 4032 47584 4060
rect 47535 4029 47547 4032
rect 47489 4023 47547 4029
rect 46477 3995 46535 4001
rect 43824 3964 45140 3992
rect 18782 3924 18788 3936
rect 16132 3896 18788 3924
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 18874 3884 18880 3936
rect 18932 3924 18938 3936
rect 20070 3924 20076 3936
rect 18932 3896 20076 3924
rect 18932 3884 18938 3896
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 20530 3924 20536 3936
rect 20491 3896 20536 3924
rect 20530 3884 20536 3896
rect 20588 3884 20594 3936
rect 22646 3924 22652 3936
rect 22607 3896 22652 3924
rect 22646 3884 22652 3896
rect 22704 3884 22710 3936
rect 27246 3924 27252 3936
rect 27207 3896 27252 3924
rect 27246 3884 27252 3896
rect 27304 3884 27310 3936
rect 27338 3884 27344 3936
rect 27396 3924 27402 3936
rect 31846 3924 31852 3936
rect 27396 3896 31852 3924
rect 27396 3884 27402 3896
rect 31846 3884 31852 3896
rect 31904 3884 31910 3936
rect 32030 3884 32036 3936
rect 32088 3924 32094 3936
rect 32674 3924 32680 3936
rect 32088 3896 32680 3924
rect 32088 3884 32094 3896
rect 32674 3884 32680 3896
rect 32732 3924 32738 3936
rect 32861 3927 32919 3933
rect 32861 3924 32873 3927
rect 32732 3896 32873 3924
rect 32732 3884 32738 3896
rect 32861 3893 32873 3896
rect 32907 3924 32919 3927
rect 34422 3924 34428 3936
rect 32907 3896 34428 3924
rect 32907 3893 32919 3896
rect 32861 3887 32919 3893
rect 34422 3884 34428 3896
rect 34480 3884 34486 3936
rect 35710 3884 35716 3936
rect 35768 3924 35774 3936
rect 36081 3927 36139 3933
rect 36081 3924 36093 3927
rect 35768 3896 36093 3924
rect 35768 3884 35774 3896
rect 36081 3893 36093 3896
rect 36127 3893 36139 3927
rect 36081 3887 36139 3893
rect 36170 3884 36176 3936
rect 36228 3924 36234 3936
rect 41138 3924 41144 3936
rect 36228 3896 41144 3924
rect 36228 3884 36234 3896
rect 41138 3884 41144 3896
rect 41196 3884 41202 3936
rect 41230 3884 41236 3936
rect 41288 3924 41294 3936
rect 45112 3933 45140 3964
rect 46477 3961 46489 3995
rect 46523 3992 46535 3995
rect 46566 3992 46572 4004
rect 46523 3964 46572 3992
rect 46523 3961 46535 3964
rect 46477 3955 46535 3961
rect 46566 3952 46572 3964
rect 46624 3952 46630 4004
rect 47136 3992 47164 4023
rect 47578 4020 47584 4032
rect 47636 4020 47642 4072
rect 47673 4063 47731 4069
rect 47673 4029 47685 4063
rect 47719 4060 47731 4063
rect 49510 4060 49516 4072
rect 47719 4032 49516 4060
rect 47719 4029 47731 4032
rect 47673 4023 47731 4029
rect 49510 4020 49516 4032
rect 49568 4020 49574 4072
rect 49620 4069 49648 4100
rect 51718 4088 51724 4140
rect 51776 4128 51782 4140
rect 52273 4131 52331 4137
rect 52273 4128 52285 4131
rect 51776 4100 52285 4128
rect 51776 4088 51782 4100
rect 52273 4097 52285 4100
rect 52319 4097 52331 4131
rect 54018 4128 54024 4140
rect 52273 4091 52331 4097
rect 52380 4100 54024 4128
rect 49605 4063 49663 4069
rect 49605 4029 49617 4063
rect 49651 4029 49663 4063
rect 49605 4023 49663 4029
rect 49789 4063 49847 4069
rect 49789 4029 49801 4063
rect 49835 4060 49847 4063
rect 49878 4060 49884 4072
rect 49835 4032 49884 4060
rect 49835 4029 49847 4032
rect 49789 4023 49847 4029
rect 49878 4020 49884 4032
rect 49936 4020 49942 4072
rect 49973 4063 50031 4069
rect 49973 4029 49985 4063
rect 50019 4060 50031 4063
rect 50062 4060 50068 4072
rect 50019 4032 50068 4060
rect 50019 4029 50031 4032
rect 49973 4023 50031 4029
rect 50062 4020 50068 4032
rect 50120 4020 50126 4072
rect 48222 3992 48228 4004
rect 47136 3964 48228 3992
rect 48222 3952 48228 3964
rect 48280 3992 48286 4004
rect 52380 3992 52408 4100
rect 54018 4088 54024 4100
rect 54076 4088 54082 4140
rect 55306 4088 55312 4140
rect 55364 4128 55370 4140
rect 55493 4131 55551 4137
rect 55493 4128 55505 4131
rect 55364 4100 55505 4128
rect 55364 4088 55370 4100
rect 55493 4097 55505 4100
rect 55539 4128 55551 4131
rect 56686 4128 56692 4140
rect 55539 4100 56692 4128
rect 55539 4097 55551 4100
rect 55493 4091 55551 4097
rect 56686 4088 56692 4100
rect 56744 4088 56750 4140
rect 59446 4128 59452 4140
rect 56796 4100 59452 4128
rect 52549 4063 52607 4069
rect 52549 4029 52561 4063
rect 52595 4060 52607 4063
rect 53466 4060 53472 4072
rect 52595 4032 53472 4060
rect 52595 4029 52607 4032
rect 52549 4023 52607 4029
rect 53466 4020 53472 4032
rect 53524 4020 53530 4072
rect 55398 4060 55404 4072
rect 55359 4032 55404 4060
rect 55398 4020 55404 4032
rect 55456 4020 55462 4072
rect 55858 4060 55864 4072
rect 55819 4032 55864 4060
rect 55858 4020 55864 4032
rect 55916 4020 55922 4072
rect 55950 4020 55956 4072
rect 56008 4060 56014 4072
rect 56796 4060 56824 4100
rect 59446 4088 59452 4100
rect 59504 4088 59510 4140
rect 56008 4032 56824 4060
rect 57425 4063 57483 4069
rect 56008 4020 56014 4032
rect 57425 4029 57437 4063
rect 57471 4060 57483 4063
rect 57790 4060 57796 4072
rect 57471 4032 57796 4060
rect 57471 4029 57483 4032
rect 57425 4023 57483 4029
rect 57790 4020 57796 4032
rect 57848 4020 57854 4072
rect 58526 4060 58532 4072
rect 58487 4032 58532 4060
rect 58526 4020 58532 4032
rect 58584 4020 58590 4072
rect 58802 4060 58808 4072
rect 58763 4032 58808 4060
rect 58802 4020 58808 4032
rect 58860 4020 58866 4072
rect 48280 3964 52408 3992
rect 53208 3964 57652 3992
rect 48280 3952 48286 3964
rect 41969 3927 42027 3933
rect 41969 3924 41981 3927
rect 41288 3896 41981 3924
rect 41288 3884 41294 3896
rect 41969 3893 41981 3896
rect 42015 3893 42027 3927
rect 41969 3887 42027 3893
rect 45097 3927 45155 3933
rect 45097 3893 45109 3927
rect 45143 3924 45155 3927
rect 45646 3924 45652 3936
rect 45143 3896 45652 3924
rect 45143 3893 45155 3896
rect 45097 3887 45155 3893
rect 45646 3884 45652 3896
rect 45704 3884 45710 3936
rect 51626 3884 51632 3936
rect 51684 3924 51690 3936
rect 53208 3924 53236 3964
rect 51684 3896 53236 3924
rect 51684 3884 51690 3896
rect 53742 3884 53748 3936
rect 53800 3924 53806 3936
rect 53837 3927 53895 3933
rect 53837 3924 53849 3927
rect 53800 3896 53849 3924
rect 53800 3884 53806 3896
rect 53837 3893 53849 3896
rect 53883 3893 53895 3927
rect 53837 3887 53895 3893
rect 55582 3884 55588 3936
rect 55640 3924 55646 3936
rect 55950 3924 55956 3936
rect 55640 3896 55956 3924
rect 55640 3884 55646 3896
rect 55950 3884 55956 3896
rect 56008 3884 56014 3936
rect 57624 3933 57652 3964
rect 57609 3927 57667 3933
rect 57609 3893 57621 3927
rect 57655 3924 57667 3927
rect 57698 3924 57704 3936
rect 57655 3896 57704 3924
rect 57655 3893 57667 3896
rect 57609 3887 57667 3893
rect 57698 3884 57704 3896
rect 57756 3884 57762 3936
rect 57974 3884 57980 3936
rect 58032 3924 58038 3936
rect 59909 3927 59967 3933
rect 59909 3924 59921 3927
rect 58032 3896 59921 3924
rect 58032 3884 58038 3896
rect 59909 3893 59921 3896
rect 59955 3893 59967 3927
rect 59909 3887 59967 3893
rect 1104 3834 62192 3856
rect 1104 3782 21344 3834
rect 21396 3782 21408 3834
rect 21460 3782 21472 3834
rect 21524 3782 21536 3834
rect 21588 3782 41707 3834
rect 41759 3782 41771 3834
rect 41823 3782 41835 3834
rect 41887 3782 41899 3834
rect 41951 3782 62192 3834
rect 1104 3760 62192 3782
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 14182 3720 14188 3732
rect 4028 3692 14188 3720
rect 4028 3680 4034 3692
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 16022 3680 16028 3732
rect 16080 3720 16086 3732
rect 19058 3720 19064 3732
rect 16080 3692 19064 3720
rect 16080 3680 16086 3692
rect 19058 3680 19064 3692
rect 19116 3720 19122 3732
rect 21082 3720 21088 3732
rect 19116 3692 21088 3720
rect 19116 3680 19122 3692
rect 21082 3680 21088 3692
rect 21140 3680 21146 3732
rect 23474 3720 23480 3732
rect 23435 3692 23480 3720
rect 23474 3680 23480 3692
rect 23532 3680 23538 3732
rect 25498 3680 25504 3732
rect 25556 3720 25562 3732
rect 27338 3720 27344 3732
rect 25556 3692 27344 3720
rect 25556 3680 25562 3692
rect 27338 3680 27344 3692
rect 27396 3680 27402 3732
rect 27798 3720 27804 3732
rect 27759 3692 27804 3720
rect 27798 3680 27804 3692
rect 27856 3680 27862 3732
rect 29564 3692 29960 3720
rect 6638 3652 6644 3664
rect 4540 3624 6644 3652
rect 4540 3593 4568 3624
rect 6638 3612 6644 3624
rect 6696 3612 6702 3664
rect 6730 3612 6736 3664
rect 6788 3652 6794 3664
rect 12710 3652 12716 3664
rect 6788 3624 12716 3652
rect 6788 3612 6794 3624
rect 12710 3612 12716 3624
rect 12768 3612 12774 3664
rect 12986 3612 12992 3664
rect 13044 3652 13050 3664
rect 22646 3652 22652 3664
rect 13044 3624 22652 3652
rect 13044 3612 13050 3624
rect 22646 3612 22652 3624
rect 22704 3652 22710 3664
rect 27706 3652 27712 3664
rect 22704 3624 25452 3652
rect 27667 3624 27712 3652
rect 22704 3612 22710 3624
rect 4525 3587 4583 3593
rect 4525 3553 4537 3587
rect 4571 3553 4583 3587
rect 6454 3584 6460 3596
rect 6415 3556 6460 3584
rect 4525 3547 4583 3553
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 6825 3587 6883 3593
rect 6825 3553 6837 3587
rect 6871 3553 6883 3587
rect 6825 3547 6883 3553
rect 7009 3587 7067 3593
rect 7009 3553 7021 3587
rect 7055 3584 7067 3587
rect 7374 3584 7380 3596
rect 7055 3556 7380 3584
rect 7055 3553 7067 3556
rect 7009 3547 7067 3553
rect 4433 3519 4491 3525
rect 4433 3485 4445 3519
rect 4479 3485 4491 3519
rect 4982 3516 4988 3528
rect 4943 3488 4988 3516
rect 4433 3479 4491 3485
rect 4448 3448 4476 3479
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 6546 3516 6552 3528
rect 6507 3488 6552 3516
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 6840 3516 6868 3547
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 7926 3584 7932 3596
rect 7887 3556 7932 3584
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 8570 3584 8576 3596
rect 8531 3556 8576 3584
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 11977 3587 12035 3593
rect 11977 3553 11989 3587
rect 12023 3584 12035 3587
rect 12802 3584 12808 3596
rect 12023 3556 12808 3584
rect 12023 3553 12035 3556
rect 11977 3547 12035 3553
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 13078 3584 13084 3596
rect 13039 3556 13084 3584
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 13265 3587 13323 3593
rect 13265 3553 13277 3587
rect 13311 3553 13323 3587
rect 16298 3584 16304 3596
rect 16259 3556 16304 3584
rect 13265 3547 13323 3553
rect 6840 3488 8064 3516
rect 8036 3460 8064 3488
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 10778 3516 10784 3528
rect 8260 3488 10784 3516
rect 8260 3476 8266 3488
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 13280 3516 13308 3547
rect 16298 3544 16304 3556
rect 16356 3544 16362 3596
rect 16485 3587 16543 3593
rect 16485 3553 16497 3587
rect 16531 3553 16543 3587
rect 16485 3547 16543 3553
rect 12492 3488 13308 3516
rect 13633 3519 13691 3525
rect 12492 3476 12498 3488
rect 13633 3485 13645 3519
rect 13679 3516 13691 3519
rect 13722 3516 13728 3528
rect 13679 3488 13728 3516
rect 13679 3485 13691 3488
rect 13633 3479 13691 3485
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 15562 3476 15568 3528
rect 15620 3516 15626 3528
rect 16500 3516 16528 3547
rect 16850 3544 16856 3596
rect 16908 3584 16914 3596
rect 17037 3587 17095 3593
rect 17037 3584 17049 3587
rect 16908 3556 17049 3584
rect 16908 3544 16914 3556
rect 17037 3553 17049 3556
rect 17083 3553 17095 3587
rect 17218 3584 17224 3596
rect 17179 3556 17224 3584
rect 17037 3547 17095 3553
rect 17218 3544 17224 3556
rect 17276 3584 17282 3596
rect 18874 3584 18880 3596
rect 17276 3556 18736 3584
rect 18835 3556 18880 3584
rect 17276 3544 17282 3556
rect 15620 3488 16528 3516
rect 15620 3476 15626 3488
rect 17494 3476 17500 3528
rect 17552 3516 17558 3528
rect 18506 3516 18512 3528
rect 17552 3488 18512 3516
rect 17552 3476 17558 3488
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 18601 3519 18659 3525
rect 18601 3485 18613 3519
rect 18647 3485 18659 3519
rect 18601 3479 18659 3485
rect 5350 3448 5356 3460
rect 4448 3420 5356 3448
rect 5350 3408 5356 3420
rect 5408 3448 5414 3460
rect 5408 3420 6040 3448
rect 5408 3408 5414 3420
rect 5534 3340 5540 3392
rect 5592 3380 5598 3392
rect 5905 3383 5963 3389
rect 5905 3380 5917 3383
rect 5592 3352 5917 3380
rect 5592 3340 5598 3352
rect 5905 3349 5917 3352
rect 5951 3349 5963 3383
rect 6012 3380 6040 3420
rect 7466 3408 7472 3460
rect 7524 3448 7530 3460
rect 7834 3448 7840 3460
rect 7524 3420 7840 3448
rect 7524 3408 7530 3420
rect 7834 3408 7840 3420
rect 7892 3448 7898 3460
rect 7929 3451 7987 3457
rect 7929 3448 7941 3451
rect 7892 3420 7941 3448
rect 7892 3408 7898 3420
rect 7929 3417 7941 3420
rect 7975 3417 7987 3451
rect 7929 3411 7987 3417
rect 8018 3408 8024 3460
rect 8076 3448 8082 3460
rect 16022 3448 16028 3460
rect 8076 3420 16028 3448
rect 8076 3408 8082 3420
rect 16022 3408 16028 3420
rect 16080 3408 16086 3460
rect 16298 3408 16304 3460
rect 16356 3448 16362 3460
rect 17770 3448 17776 3460
rect 16356 3420 17776 3448
rect 16356 3408 16362 3420
rect 17770 3408 17776 3420
rect 17828 3408 17834 3460
rect 18230 3408 18236 3460
rect 18288 3448 18294 3460
rect 18616 3448 18644 3479
rect 18288 3420 18644 3448
rect 18708 3448 18736 3556
rect 18874 3544 18880 3556
rect 18932 3584 18938 3596
rect 19242 3584 19248 3596
rect 18932 3556 19248 3584
rect 18932 3544 18938 3556
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 19334 3544 19340 3596
rect 19392 3584 19398 3596
rect 20898 3584 20904 3596
rect 19392 3556 19437 3584
rect 20859 3556 20904 3584
rect 19392 3544 19398 3556
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 23198 3584 23204 3596
rect 23159 3556 23204 3584
rect 23198 3544 23204 3556
rect 23256 3544 23262 3596
rect 23385 3587 23443 3593
rect 23385 3553 23397 3587
rect 23431 3584 23443 3587
rect 24210 3584 24216 3596
rect 23431 3556 24216 3584
rect 23431 3553 23443 3556
rect 23385 3547 23443 3553
rect 19613 3519 19671 3525
rect 19613 3485 19625 3519
rect 19659 3516 19671 3519
rect 20714 3516 20720 3528
rect 19659 3488 20720 3516
rect 19659 3485 19671 3488
rect 19613 3479 19671 3485
rect 20714 3476 20720 3488
rect 20772 3476 20778 3528
rect 22830 3476 22836 3528
rect 22888 3516 22894 3528
rect 23400 3516 23428 3547
rect 24210 3544 24216 3556
rect 24268 3544 24274 3596
rect 25424 3593 25452 3624
rect 27706 3612 27712 3624
rect 27764 3612 27770 3664
rect 27890 3652 27896 3664
rect 27851 3624 27896 3652
rect 27890 3612 27896 3624
rect 27948 3612 27954 3664
rect 28258 3652 28264 3664
rect 28219 3624 28264 3652
rect 28258 3612 28264 3624
rect 28316 3612 28322 3664
rect 25409 3587 25467 3593
rect 25409 3553 25421 3587
rect 25455 3553 25467 3587
rect 25409 3547 25467 3553
rect 22888 3488 23428 3516
rect 24581 3519 24639 3525
rect 22888 3476 22894 3488
rect 24581 3485 24593 3519
rect 24627 3516 24639 3519
rect 24854 3516 24860 3528
rect 24627 3488 24860 3516
rect 24627 3485 24639 3488
rect 24581 3479 24639 3485
rect 24854 3476 24860 3488
rect 24912 3476 24918 3528
rect 25133 3519 25191 3525
rect 25133 3485 25145 3519
rect 25179 3485 25191 3519
rect 25133 3479 25191 3485
rect 25593 3519 25651 3525
rect 25593 3485 25605 3519
rect 25639 3516 25651 3519
rect 26234 3516 26240 3528
rect 25639 3488 26240 3516
rect 25639 3485 25651 3488
rect 25593 3479 25651 3485
rect 20622 3448 20628 3460
rect 18708 3420 20628 3448
rect 18288 3408 18294 3420
rect 9122 3380 9128 3392
rect 6012 3352 9128 3380
rect 5905 3343 5963 3349
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 12161 3383 12219 3389
rect 12161 3349 12173 3383
rect 12207 3380 12219 3383
rect 13262 3380 13268 3392
rect 12207 3352 13268 3380
rect 12207 3349 12219 3352
rect 12161 3343 12219 3349
rect 13262 3340 13268 3352
rect 13320 3340 13326 3392
rect 13906 3340 13912 3392
rect 13964 3380 13970 3392
rect 17497 3383 17555 3389
rect 17497 3380 17509 3383
rect 13964 3352 17509 3380
rect 13964 3340 13970 3352
rect 17497 3349 17509 3352
rect 17543 3349 17555 3383
rect 18616 3380 18644 3420
rect 20622 3408 20628 3420
rect 20680 3408 20686 3460
rect 25148 3448 25176 3479
rect 26234 3476 26240 3488
rect 26292 3476 26298 3528
rect 27522 3516 27528 3528
rect 27483 3488 27528 3516
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 27724 3516 27752 3612
rect 29564 3516 29592 3692
rect 29730 3612 29736 3664
rect 29788 3652 29794 3664
rect 29825 3655 29883 3661
rect 29825 3652 29837 3655
rect 29788 3624 29837 3652
rect 29788 3612 29794 3624
rect 29825 3621 29837 3624
rect 29871 3621 29883 3655
rect 29932 3652 29960 3692
rect 30098 3680 30104 3732
rect 30156 3720 30162 3732
rect 32217 3723 32275 3729
rect 32217 3720 32229 3723
rect 30156 3692 32229 3720
rect 30156 3680 30162 3692
rect 32217 3689 32229 3692
rect 32263 3689 32275 3723
rect 34333 3723 34391 3729
rect 34333 3720 34345 3723
rect 32217 3683 32275 3689
rect 32784 3692 34345 3720
rect 29932 3624 32720 3652
rect 29825 3615 29883 3621
rect 29917 3587 29975 3593
rect 29917 3553 29929 3587
rect 29963 3584 29975 3587
rect 30006 3584 30012 3596
rect 29963 3556 30012 3584
rect 29963 3553 29975 3556
rect 29917 3547 29975 3553
rect 30006 3544 30012 3556
rect 30064 3544 30070 3596
rect 27724 3488 29592 3516
rect 29641 3519 29699 3525
rect 29641 3485 29653 3519
rect 29687 3516 29699 3519
rect 31110 3516 31116 3528
rect 29687 3488 31116 3516
rect 29687 3485 29699 3488
rect 29641 3479 29699 3485
rect 31110 3476 31116 3488
rect 31168 3476 31174 3528
rect 32306 3476 32312 3528
rect 32364 3516 32370 3528
rect 32585 3519 32643 3525
rect 32585 3516 32597 3519
rect 32364 3488 32597 3516
rect 32364 3476 32370 3488
rect 32585 3485 32597 3488
rect 32631 3485 32643 3519
rect 32692 3516 32720 3624
rect 32784 3593 32812 3692
rect 34333 3689 34345 3692
rect 34379 3720 34391 3723
rect 39574 3720 39580 3732
rect 34379 3692 39580 3720
rect 34379 3689 34391 3692
rect 34333 3683 34391 3689
rect 39574 3680 39580 3692
rect 39632 3720 39638 3732
rect 40313 3723 40371 3729
rect 40313 3720 40325 3723
rect 39632 3692 40325 3720
rect 39632 3680 39638 3692
rect 40313 3689 40325 3692
rect 40359 3689 40371 3723
rect 41598 3720 41604 3732
rect 41559 3692 41604 3720
rect 40313 3683 40371 3689
rect 41598 3680 41604 3692
rect 41656 3680 41662 3732
rect 43346 3680 43352 3732
rect 43404 3720 43410 3732
rect 49694 3720 49700 3732
rect 43404 3692 49700 3720
rect 43404 3680 43410 3692
rect 49694 3680 49700 3692
rect 49752 3680 49758 3732
rect 49878 3720 49884 3732
rect 49839 3692 49884 3720
rect 49878 3680 49884 3692
rect 49936 3680 49942 3732
rect 57606 3680 57612 3732
rect 57664 3720 57670 3732
rect 57664 3692 59216 3720
rect 57664 3680 57670 3692
rect 34517 3655 34575 3661
rect 34517 3652 34529 3655
rect 33244 3624 34529 3652
rect 32769 3587 32827 3593
rect 32769 3553 32781 3587
rect 32815 3553 32827 3587
rect 33137 3587 33195 3593
rect 33137 3584 33149 3587
rect 32769 3547 32827 3553
rect 32876 3556 33149 3584
rect 32876 3516 32904 3556
rect 33137 3553 33149 3556
rect 33183 3553 33195 3587
rect 33137 3547 33195 3553
rect 33042 3516 33048 3528
rect 32692 3488 32904 3516
rect 33003 3488 33048 3516
rect 32585 3479 32643 3485
rect 33042 3476 33048 3488
rect 33100 3516 33106 3528
rect 33244 3516 33272 3624
rect 34517 3621 34529 3624
rect 34563 3621 34575 3655
rect 34517 3615 34575 3621
rect 34606 3612 34612 3664
rect 34664 3652 34670 3664
rect 34885 3655 34943 3661
rect 34885 3652 34897 3655
rect 34664 3624 34897 3652
rect 34664 3612 34670 3624
rect 34885 3621 34897 3624
rect 34931 3621 34943 3655
rect 35989 3655 36047 3661
rect 35989 3652 36001 3655
rect 34885 3615 34943 3621
rect 35544 3624 36001 3652
rect 34422 3584 34428 3596
rect 33100 3488 33272 3516
rect 34072 3556 34284 3584
rect 34383 3556 34428 3584
rect 33100 3476 33106 3488
rect 30558 3448 30564 3460
rect 25148 3420 30564 3448
rect 30558 3408 30564 3420
rect 30616 3408 30622 3460
rect 30742 3408 30748 3460
rect 30800 3448 30806 3460
rect 34072 3448 34100 3556
rect 34149 3519 34207 3525
rect 34149 3485 34161 3519
rect 34195 3485 34207 3519
rect 34149 3479 34207 3485
rect 30800 3420 34100 3448
rect 30800 3408 30806 3420
rect 19702 3380 19708 3392
rect 18616 3352 19708 3380
rect 17497 3343 17555 3349
rect 19702 3340 19708 3352
rect 19760 3380 19766 3392
rect 20346 3380 20352 3392
rect 19760 3352 20352 3380
rect 19760 3340 19766 3352
rect 20346 3340 20352 3352
rect 20404 3340 20410 3392
rect 22462 3340 22468 3392
rect 22520 3380 22526 3392
rect 29270 3380 29276 3392
rect 22520 3352 29276 3380
rect 22520 3340 22526 3352
rect 29270 3340 29276 3352
rect 29328 3340 29334 3392
rect 29362 3340 29368 3392
rect 29420 3380 29426 3392
rect 30101 3383 30159 3389
rect 30101 3380 30113 3383
rect 29420 3352 30113 3380
rect 29420 3340 29426 3352
rect 30101 3349 30113 3352
rect 30147 3349 30159 3383
rect 30101 3343 30159 3349
rect 31294 3340 31300 3392
rect 31352 3380 31358 3392
rect 32398 3380 32404 3392
rect 31352 3352 32404 3380
rect 31352 3340 31358 3352
rect 32398 3340 32404 3352
rect 32456 3340 32462 3392
rect 32950 3340 32956 3392
rect 33008 3380 33014 3392
rect 34164 3380 34192 3479
rect 34256 3448 34284 3556
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 35544 3528 35572 3624
rect 35989 3621 36001 3624
rect 36035 3621 36047 3655
rect 35989 3615 36047 3621
rect 36081 3655 36139 3661
rect 36081 3621 36093 3655
rect 36127 3652 36139 3655
rect 36170 3652 36176 3664
rect 36127 3624 36176 3652
rect 36127 3621 36139 3624
rect 36081 3615 36139 3621
rect 36170 3612 36176 3624
rect 36228 3612 36234 3664
rect 36262 3612 36268 3664
rect 36320 3652 36326 3664
rect 38838 3652 38844 3664
rect 36320 3624 38844 3652
rect 36320 3612 36326 3624
rect 38838 3612 38844 3624
rect 38896 3612 38902 3664
rect 52917 3655 52975 3661
rect 52917 3621 52929 3655
rect 52963 3652 52975 3655
rect 55858 3652 55864 3664
rect 52963 3624 55864 3652
rect 52963 3621 52975 3624
rect 52917 3615 52975 3621
rect 55858 3612 55864 3624
rect 55916 3612 55922 3664
rect 58069 3655 58127 3661
rect 58069 3621 58081 3655
rect 58115 3652 58127 3655
rect 58802 3652 58808 3664
rect 58115 3624 58808 3652
rect 58115 3621 58127 3624
rect 58069 3615 58127 3621
rect 58802 3612 58808 3624
rect 58860 3612 58866 3664
rect 35897 3587 35955 3593
rect 35897 3553 35909 3587
rect 35943 3584 35955 3587
rect 35943 3556 36676 3584
rect 35943 3553 35955 3556
rect 35897 3547 35955 3553
rect 35526 3516 35532 3528
rect 35487 3488 35532 3516
rect 35526 3476 35532 3488
rect 35584 3476 35590 3528
rect 35713 3519 35771 3525
rect 35713 3485 35725 3519
rect 35759 3516 35771 3519
rect 36354 3516 36360 3528
rect 35759 3488 36360 3516
rect 35759 3485 35771 3488
rect 35713 3479 35771 3485
rect 36354 3476 36360 3488
rect 36412 3476 36418 3528
rect 36449 3519 36507 3525
rect 36449 3485 36461 3519
rect 36495 3485 36507 3519
rect 36648 3516 36676 3556
rect 36722 3544 36728 3596
rect 36780 3584 36786 3596
rect 37182 3584 37188 3596
rect 36780 3556 37188 3584
rect 36780 3544 36786 3556
rect 37182 3544 37188 3556
rect 37240 3584 37246 3596
rect 37737 3587 37795 3593
rect 37737 3584 37749 3587
rect 37240 3556 37749 3584
rect 37240 3544 37246 3556
rect 37737 3553 37749 3556
rect 37783 3553 37795 3587
rect 37737 3547 37795 3553
rect 37826 3544 37832 3596
rect 37884 3584 37890 3596
rect 39022 3584 39028 3596
rect 37884 3556 39028 3584
rect 37884 3544 37890 3556
rect 39022 3544 39028 3556
rect 39080 3544 39086 3596
rect 39206 3584 39212 3596
rect 39167 3556 39212 3584
rect 39206 3544 39212 3556
rect 39264 3544 39270 3596
rect 40402 3544 40408 3596
rect 40460 3584 40466 3596
rect 41417 3587 41475 3593
rect 41417 3584 41429 3587
rect 40460 3556 41429 3584
rect 40460 3544 40466 3556
rect 41417 3553 41429 3556
rect 41463 3553 41475 3587
rect 41417 3547 41475 3553
rect 43622 3544 43628 3596
rect 43680 3584 43686 3596
rect 44082 3584 44088 3596
rect 43680 3556 44088 3584
rect 43680 3544 43686 3556
rect 44082 3544 44088 3556
rect 44140 3584 44146 3596
rect 45189 3587 45247 3593
rect 45189 3584 45201 3587
rect 44140 3556 45201 3584
rect 44140 3544 44146 3556
rect 45189 3553 45201 3556
rect 45235 3553 45247 3587
rect 46566 3584 46572 3596
rect 46527 3556 46572 3584
rect 45189 3547 45247 3553
rect 46566 3544 46572 3556
rect 46624 3544 46630 3596
rect 49605 3587 49663 3593
rect 49605 3553 49617 3587
rect 49651 3553 49663 3587
rect 49605 3547 49663 3553
rect 38470 3516 38476 3528
rect 36648 3488 38476 3516
rect 36449 3479 36507 3485
rect 36464 3448 36492 3479
rect 38470 3476 38476 3488
rect 38528 3476 38534 3528
rect 38933 3519 38991 3525
rect 38933 3485 38945 3519
rect 38979 3485 38991 3519
rect 38933 3479 38991 3485
rect 34256 3420 36492 3448
rect 36556 3420 38056 3448
rect 36556 3380 36584 3420
rect 33008 3352 36584 3380
rect 33008 3340 33014 3352
rect 37642 3340 37648 3392
rect 37700 3380 37706 3392
rect 37921 3383 37979 3389
rect 37921 3380 37933 3383
rect 37700 3352 37933 3380
rect 37700 3340 37706 3352
rect 37921 3349 37933 3352
rect 37967 3349 37979 3383
rect 38028 3380 38056 3420
rect 38562 3408 38568 3460
rect 38620 3448 38626 3460
rect 38948 3448 38976 3479
rect 40494 3476 40500 3528
rect 40552 3516 40558 3528
rect 46106 3516 46112 3528
rect 40552 3488 46112 3516
rect 40552 3476 40558 3488
rect 46106 3476 46112 3488
rect 46164 3516 46170 3528
rect 46293 3519 46351 3525
rect 46293 3516 46305 3519
rect 46164 3488 46305 3516
rect 46164 3476 46170 3488
rect 46293 3485 46305 3488
rect 46339 3485 46351 3519
rect 49620 3516 49648 3547
rect 49694 3544 49700 3596
rect 49752 3584 49758 3596
rect 49789 3587 49847 3593
rect 49789 3584 49801 3587
rect 49752 3556 49801 3584
rect 49752 3544 49758 3556
rect 49789 3553 49801 3556
rect 49835 3584 49847 3587
rect 51626 3584 51632 3596
rect 49835 3556 51632 3584
rect 49835 3553 49847 3556
rect 49789 3547 49847 3553
rect 51626 3544 51632 3556
rect 51684 3544 51690 3596
rect 55306 3584 55312 3596
rect 55267 3556 55312 3584
rect 55306 3544 55312 3556
rect 55364 3544 55370 3596
rect 55674 3584 55680 3596
rect 55635 3556 55680 3584
rect 55674 3544 55680 3556
rect 55732 3544 55738 3596
rect 56778 3584 56784 3596
rect 56739 3556 56784 3584
rect 56778 3544 56784 3556
rect 56836 3544 56842 3596
rect 56870 3544 56876 3596
rect 56928 3584 56934 3596
rect 58710 3584 58716 3596
rect 56928 3556 58716 3584
rect 56928 3544 56934 3556
rect 58710 3544 58716 3556
rect 58768 3544 58774 3596
rect 58894 3544 58900 3596
rect 58952 3584 58958 3596
rect 59188 3593 59216 3692
rect 59081 3587 59139 3593
rect 59081 3584 59093 3587
rect 58952 3556 59093 3584
rect 58952 3544 58958 3556
rect 59081 3553 59093 3556
rect 59127 3553 59139 3587
rect 59081 3547 59139 3553
rect 59173 3587 59231 3593
rect 59173 3553 59185 3587
rect 59219 3553 59231 3587
rect 59173 3547 59231 3553
rect 60185 3587 60243 3593
rect 60185 3553 60197 3587
rect 60231 3584 60243 3587
rect 61010 3584 61016 3596
rect 60231 3556 61016 3584
rect 60231 3553 60243 3556
rect 60185 3547 60243 3553
rect 61010 3544 61016 3556
rect 61068 3544 61074 3596
rect 50430 3516 50436 3528
rect 49620 3488 50436 3516
rect 46293 3479 46351 3485
rect 50430 3476 50436 3488
rect 50488 3476 50494 3528
rect 51258 3476 51264 3528
rect 51316 3516 51322 3528
rect 51537 3519 51595 3525
rect 51537 3516 51549 3519
rect 51316 3488 51549 3516
rect 51316 3476 51322 3488
rect 51537 3485 51549 3488
rect 51583 3485 51595 3519
rect 51537 3479 51595 3485
rect 52089 3519 52147 3525
rect 52089 3485 52101 3519
rect 52135 3516 52147 3519
rect 52178 3516 52184 3528
rect 52135 3488 52184 3516
rect 52135 3485 52147 3488
rect 52089 3479 52147 3485
rect 52178 3476 52184 3488
rect 52236 3476 52242 3528
rect 53064 3519 53122 3525
rect 53064 3485 53076 3519
rect 53110 3516 53122 3519
rect 53190 3516 53196 3528
rect 53110 3488 53196 3516
rect 53110 3485 53122 3488
rect 53064 3479 53122 3485
rect 53190 3476 53196 3488
rect 53248 3476 53254 3528
rect 53285 3519 53343 3525
rect 53285 3485 53297 3519
rect 53331 3485 53343 3519
rect 53285 3479 53343 3485
rect 38620 3420 38976 3448
rect 38620 3408 38626 3420
rect 41138 3408 41144 3460
rect 41196 3448 41202 3460
rect 43806 3448 43812 3460
rect 41196 3420 43812 3448
rect 41196 3408 41202 3420
rect 43806 3408 43812 3420
rect 43864 3448 43870 3460
rect 45373 3451 45431 3457
rect 45373 3448 45385 3451
rect 43864 3420 45385 3448
rect 43864 3408 43870 3420
rect 45373 3417 45385 3420
rect 45419 3417 45431 3451
rect 45373 3411 45431 3417
rect 50614 3408 50620 3460
rect 50672 3448 50678 3460
rect 53300 3448 53328 3479
rect 54570 3476 54576 3528
rect 54628 3516 54634 3528
rect 54665 3519 54723 3525
rect 54665 3516 54677 3519
rect 54628 3488 54677 3516
rect 54628 3476 54634 3488
rect 54665 3485 54677 3488
rect 54711 3485 54723 3519
rect 54665 3479 54723 3485
rect 55401 3519 55459 3525
rect 55401 3485 55413 3519
rect 55447 3485 55459 3519
rect 55582 3516 55588 3528
rect 55543 3488 55588 3516
rect 55401 3479 55459 3485
rect 50672 3420 53328 3448
rect 55416 3448 55444 3479
rect 55582 3476 55588 3488
rect 55640 3476 55646 3528
rect 55766 3476 55772 3528
rect 55824 3516 55830 3528
rect 56689 3519 56747 3525
rect 56689 3516 56701 3519
rect 55824 3488 56701 3516
rect 55824 3476 55830 3488
rect 56689 3485 56701 3488
rect 56735 3485 56747 3519
rect 56689 3479 56747 3485
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 58621 3519 58679 3525
rect 58621 3516 58633 3519
rect 58492 3488 58633 3516
rect 58492 3476 58498 3488
rect 58621 3485 58633 3488
rect 58667 3485 58679 3519
rect 58621 3479 58679 3485
rect 55416 3420 56732 3448
rect 50672 3408 50678 3420
rect 41230 3380 41236 3392
rect 38028 3352 41236 3380
rect 37921 3343 37979 3349
rect 41230 3340 41236 3352
rect 41288 3340 41294 3392
rect 47857 3383 47915 3389
rect 47857 3349 47869 3383
rect 47903 3380 47915 3383
rect 49970 3380 49976 3392
rect 47903 3352 49976 3380
rect 47903 3349 47915 3352
rect 47857 3343 47915 3349
rect 49970 3340 49976 3352
rect 50028 3340 50034 3392
rect 51534 3340 51540 3392
rect 51592 3380 51598 3392
rect 53193 3383 53251 3389
rect 53193 3380 53205 3383
rect 51592 3352 53205 3380
rect 51592 3340 51598 3352
rect 53193 3349 53205 3352
rect 53239 3349 53251 3383
rect 53558 3380 53564 3392
rect 53519 3352 53564 3380
rect 53193 3343 53251 3349
rect 53558 3340 53564 3352
rect 53616 3340 53622 3392
rect 56704 3380 56732 3420
rect 56965 3383 57023 3389
rect 56965 3380 56977 3383
rect 56704 3352 56977 3380
rect 56965 3349 56977 3352
rect 57011 3349 57023 3383
rect 56965 3343 57023 3349
rect 58710 3340 58716 3392
rect 58768 3380 58774 3392
rect 60277 3383 60335 3389
rect 60277 3380 60289 3383
rect 58768 3352 60289 3380
rect 58768 3340 58774 3352
rect 60277 3349 60289 3352
rect 60323 3349 60335 3383
rect 60277 3343 60335 3349
rect 1104 3290 62192 3312
rect 1104 3238 11163 3290
rect 11215 3238 11227 3290
rect 11279 3238 11291 3290
rect 11343 3238 11355 3290
rect 11407 3238 31526 3290
rect 31578 3238 31590 3290
rect 31642 3238 31654 3290
rect 31706 3238 31718 3290
rect 31770 3238 51888 3290
rect 51940 3238 51952 3290
rect 52004 3238 52016 3290
rect 52068 3238 52080 3290
rect 52132 3238 62192 3290
rect 1104 3216 62192 3238
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 6512 3148 7236 3176
rect 6512 3136 6518 3148
rect 6472 3108 6500 3136
rect 5368 3080 6500 3108
rect 4982 3000 4988 3052
rect 5040 3040 5046 3052
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 5040 3012 5273 3040
rect 5040 3000 5046 3012
rect 5261 3009 5273 3012
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 5368 2981 5396 3080
rect 6546 3068 6552 3120
rect 6604 3108 6610 3120
rect 7101 3111 7159 3117
rect 7101 3108 7113 3111
rect 6604 3080 7113 3108
rect 6604 3068 6610 3080
rect 7101 3077 7113 3080
rect 7147 3077 7159 3111
rect 7208 3108 7236 3148
rect 7558 3136 7564 3188
rect 7616 3176 7622 3188
rect 12986 3176 12992 3188
rect 7616 3148 12992 3176
rect 7616 3136 7622 3148
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 13136 3148 17724 3176
rect 13136 3136 13142 3148
rect 7208 3080 13124 3108
rect 7101 3071 7159 3077
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 6914 3040 6920 3052
rect 5859 3012 6920 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 6914 3000 6920 3012
rect 6972 3000 6978 3052
rect 7834 3040 7840 3052
rect 7795 3012 7840 3040
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 9858 3040 9864 3052
rect 8260 3012 9864 3040
rect 8260 3000 8266 3012
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 13096 3040 13124 3080
rect 13170 3068 13176 3120
rect 13228 3108 13234 3120
rect 14921 3111 14979 3117
rect 14921 3108 14933 3111
rect 13228 3080 14933 3108
rect 13228 3068 13234 3080
rect 14921 3077 14933 3080
rect 14967 3077 14979 3111
rect 14921 3071 14979 3077
rect 16025 3111 16083 3117
rect 16025 3077 16037 3111
rect 16071 3108 16083 3111
rect 17586 3108 17592 3120
rect 16071 3080 17592 3108
rect 16071 3077 16083 3080
rect 16025 3071 16083 3077
rect 17586 3068 17592 3080
rect 17644 3068 17650 3120
rect 17696 3108 17724 3148
rect 17770 3136 17776 3188
rect 17828 3176 17834 3188
rect 17828 3148 21128 3176
rect 17828 3136 17834 3148
rect 21100 3108 21128 3148
rect 21174 3136 21180 3188
rect 21232 3176 21238 3188
rect 22462 3176 22468 3188
rect 21232 3148 22468 3176
rect 21232 3136 21238 3148
rect 22462 3136 22468 3148
rect 22520 3136 22526 3188
rect 22649 3179 22707 3185
rect 22649 3145 22661 3179
rect 22695 3176 22707 3179
rect 23658 3176 23664 3188
rect 22695 3148 23664 3176
rect 22695 3145 22707 3148
rect 22649 3139 22707 3145
rect 23658 3136 23664 3148
rect 23716 3136 23722 3188
rect 26050 3136 26056 3188
rect 26108 3176 26114 3188
rect 27617 3179 27675 3185
rect 27617 3176 27629 3179
rect 26108 3148 27629 3176
rect 26108 3136 26114 3148
rect 27617 3145 27629 3148
rect 27663 3145 27675 3179
rect 27617 3139 27675 3145
rect 28074 3136 28080 3188
rect 28132 3176 28138 3188
rect 33226 3176 33232 3188
rect 28132 3148 33232 3176
rect 28132 3136 28138 3148
rect 33226 3136 33232 3148
rect 33284 3136 33290 3188
rect 33318 3136 33324 3188
rect 33376 3176 33382 3188
rect 33376 3148 37964 3176
rect 33376 3136 33382 3148
rect 24118 3108 24124 3120
rect 17696 3080 21036 3108
rect 21100 3080 24124 3108
rect 13096 3012 13400 3040
rect 5353 2975 5411 2981
rect 5353 2941 5365 2975
rect 5399 2941 5411 2975
rect 5353 2935 5411 2941
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 5767 2944 6776 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 4709 2907 4767 2913
rect 4709 2873 4721 2907
rect 4755 2904 4767 2907
rect 5902 2904 5908 2916
rect 4755 2876 5908 2904
rect 4755 2873 4767 2876
rect 4709 2867 4767 2873
rect 5902 2864 5908 2876
rect 5960 2864 5966 2916
rect 6748 2904 6776 2944
rect 6822 2932 6828 2984
rect 6880 2972 6886 2984
rect 7745 2975 7803 2981
rect 6880 2944 6925 2972
rect 6880 2932 6886 2944
rect 7745 2941 7757 2975
rect 7791 2972 7803 2975
rect 8018 2972 8024 2984
rect 7791 2944 8024 2972
rect 7791 2941 7803 2944
rect 7745 2935 7803 2941
rect 7760 2904 7788 2935
rect 8018 2932 8024 2944
rect 8076 2932 8082 2984
rect 8110 2932 8116 2984
rect 8168 2972 8174 2984
rect 13372 2981 13400 3012
rect 13446 3000 13452 3052
rect 13504 3040 13510 3052
rect 16577 3043 16635 3049
rect 13504 3012 13549 3040
rect 13648 3012 15332 3040
rect 13504 3000 13510 3012
rect 13357 2975 13415 2981
rect 8168 2944 13308 2972
rect 8168 2932 8174 2944
rect 6748 2876 7788 2904
rect 12713 2907 12771 2913
rect 12713 2873 12725 2907
rect 12759 2904 12771 2907
rect 12894 2904 12900 2916
rect 12759 2876 12900 2904
rect 12759 2873 12771 2876
rect 12713 2867 12771 2873
rect 12894 2864 12900 2876
rect 12952 2864 12958 2916
rect 13280 2904 13308 2944
rect 13357 2941 13369 2975
rect 13403 2972 13415 2975
rect 13648 2972 13676 3012
rect 13403 2944 13676 2972
rect 13403 2941 13415 2944
rect 13357 2935 13415 2941
rect 13722 2932 13728 2984
rect 13780 2972 13786 2984
rect 13906 2972 13912 2984
rect 13780 2944 13825 2972
rect 13867 2944 13912 2972
rect 13780 2932 13786 2944
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 14734 2972 14740 2984
rect 14695 2944 14740 2972
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 15304 2972 15332 3012
rect 16577 3009 16589 3043
rect 16623 3040 16635 3043
rect 18230 3040 18236 3052
rect 16623 3012 16896 3040
rect 16623 3009 16635 3012
rect 16577 3003 16635 3009
rect 16499 2975 16557 2981
rect 16499 2972 16511 2975
rect 15304 2944 16511 2972
rect 16499 2941 16511 2944
rect 16545 2972 16557 2975
rect 16758 2972 16764 2984
rect 16545 2944 16764 2972
rect 16545 2941 16557 2944
rect 16499 2935 16557 2941
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 13280 2876 16620 2904
rect 16592 2848 16620 2876
rect 7282 2796 7288 2848
rect 7340 2836 7346 2848
rect 16298 2836 16304 2848
rect 7340 2808 16304 2836
rect 7340 2796 7346 2808
rect 16298 2796 16304 2808
rect 16356 2796 16362 2848
rect 16574 2796 16580 2848
rect 16632 2796 16638 2848
rect 16868 2836 16896 3012
rect 16960 3012 18236 3040
rect 16960 2984 16988 3012
rect 18230 3000 18236 3012
rect 18288 3000 18294 3052
rect 18322 3000 18328 3052
rect 18380 3040 18386 3052
rect 19153 3043 19211 3049
rect 19153 3040 19165 3043
rect 18380 3012 19165 3040
rect 18380 3000 18386 3012
rect 19153 3009 19165 3012
rect 19199 3009 19211 3043
rect 21008 3040 21036 3080
rect 24118 3068 24124 3080
rect 24176 3068 24182 3120
rect 27522 3068 27528 3120
rect 27580 3108 27586 3120
rect 34882 3108 34888 3120
rect 27580 3080 34888 3108
rect 27580 3068 27586 3080
rect 21818 3040 21824 3052
rect 21008 3012 21824 3040
rect 19153 3003 19211 3009
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 24854 3040 24860 3052
rect 24815 3012 24860 3040
rect 24854 3000 24860 3012
rect 24912 3000 24918 3052
rect 16942 2932 16948 2984
rect 17000 2972 17006 2984
rect 17129 2975 17187 2981
rect 17000 2944 17045 2972
rect 17000 2932 17006 2944
rect 17129 2941 17141 2975
rect 17175 2972 17187 2975
rect 18690 2972 18696 2984
rect 17175 2944 18552 2972
rect 18651 2944 18696 2972
rect 17175 2941 17187 2944
rect 17129 2935 17187 2941
rect 17310 2864 17316 2916
rect 17368 2904 17374 2916
rect 18049 2907 18107 2913
rect 18049 2904 18061 2907
rect 17368 2876 18061 2904
rect 17368 2864 17374 2876
rect 18049 2873 18061 2876
rect 18095 2873 18107 2907
rect 18524 2904 18552 2944
rect 18690 2932 18696 2944
rect 18748 2932 18754 2984
rect 18782 2932 18788 2984
rect 18840 2972 18846 2984
rect 19058 2972 19064 2984
rect 18840 2944 18885 2972
rect 19019 2944 19064 2972
rect 18840 2932 18846 2944
rect 19058 2932 19064 2944
rect 19116 2932 19122 2984
rect 19242 2932 19248 2984
rect 19300 2972 19306 2984
rect 20533 2975 20591 2981
rect 19300 2944 20208 2972
rect 19300 2932 19306 2944
rect 20073 2907 20131 2913
rect 20073 2904 20085 2907
rect 18524 2876 20085 2904
rect 18049 2867 18107 2873
rect 20073 2873 20085 2876
rect 20119 2873 20131 2907
rect 20180 2904 20208 2944
rect 20533 2941 20545 2975
rect 20579 2972 20591 2975
rect 20622 2972 20628 2984
rect 20579 2944 20628 2972
rect 20579 2941 20591 2944
rect 20533 2935 20591 2941
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 20717 2975 20775 2981
rect 20717 2941 20729 2975
rect 20763 2941 20775 2975
rect 20717 2935 20775 2941
rect 20732 2904 20760 2935
rect 20806 2932 20812 2984
rect 20864 2972 20870 2984
rect 20901 2975 20959 2981
rect 20901 2972 20913 2975
rect 20864 2944 20913 2972
rect 20864 2932 20870 2944
rect 20901 2941 20913 2944
rect 20947 2941 20959 2975
rect 20901 2935 20959 2941
rect 22465 2975 22523 2981
rect 22465 2941 22477 2975
rect 22511 2972 22523 2975
rect 22554 2972 22560 2984
rect 22511 2944 22560 2972
rect 22511 2941 22523 2944
rect 22465 2935 22523 2941
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 24302 2932 24308 2984
rect 24360 2972 24366 2984
rect 27816 2981 27844 3080
rect 34882 3068 34888 3080
rect 34940 3108 34946 3120
rect 35986 3108 35992 3120
rect 34940 3080 35992 3108
rect 34940 3068 34946 3080
rect 35986 3068 35992 3080
rect 36044 3068 36050 3120
rect 36630 3108 36636 3120
rect 36096 3080 36636 3108
rect 28350 3040 28356 3052
rect 28311 3012 28356 3040
rect 28350 3000 28356 3012
rect 28408 3000 28414 3052
rect 28994 3000 29000 3052
rect 29052 3040 29058 3052
rect 30282 3040 30288 3052
rect 29052 3012 30288 3040
rect 29052 3000 29058 3012
rect 30282 3000 30288 3012
rect 30340 3000 30346 3052
rect 30466 3040 30472 3052
rect 30427 3012 30472 3040
rect 30466 3000 30472 3012
rect 30524 3000 30530 3052
rect 30926 3040 30932 3052
rect 30887 3012 30932 3040
rect 30926 3000 30932 3012
rect 30984 3000 30990 3052
rect 31018 3000 31024 3052
rect 31076 3040 31082 3052
rect 31757 3043 31815 3049
rect 31757 3040 31769 3043
rect 31076 3012 31769 3040
rect 31076 3000 31082 3012
rect 31757 3009 31769 3012
rect 31803 3009 31815 3043
rect 31757 3003 31815 3009
rect 32122 3000 32128 3052
rect 32180 3040 32186 3052
rect 32217 3043 32275 3049
rect 32217 3040 32229 3043
rect 32180 3012 32229 3040
rect 32180 3000 32186 3012
rect 32217 3009 32229 3012
rect 32263 3009 32275 3043
rect 34330 3040 34336 3052
rect 32217 3003 32275 3009
rect 32324 3012 34336 3040
rect 24581 2975 24639 2981
rect 24581 2972 24593 2975
rect 24360 2944 24593 2972
rect 24360 2932 24366 2944
rect 24581 2941 24593 2944
rect 24627 2941 24639 2975
rect 24581 2935 24639 2941
rect 27801 2975 27859 2981
rect 27801 2941 27813 2975
rect 27847 2941 27859 2975
rect 27801 2935 27859 2941
rect 27890 2932 27896 2984
rect 27948 2972 27954 2984
rect 30006 2972 30012 2984
rect 27948 2944 30012 2972
rect 27948 2932 27954 2944
rect 30006 2932 30012 2944
rect 30064 2932 30070 2984
rect 30742 2972 30748 2984
rect 30703 2944 30748 2972
rect 30742 2932 30748 2944
rect 30800 2932 30806 2984
rect 32324 2972 32352 3012
rect 30852 2944 32352 2972
rect 32401 2975 32459 2981
rect 26234 2904 26240 2916
rect 20180 2876 20760 2904
rect 26147 2876 26240 2904
rect 20073 2867 20131 2873
rect 26234 2864 26240 2876
rect 26292 2904 26298 2916
rect 29917 2907 29975 2913
rect 26292 2876 28304 2904
rect 26292 2864 26298 2876
rect 17954 2836 17960 2848
rect 16868 2808 17960 2836
rect 17954 2796 17960 2808
rect 18012 2796 18018 2848
rect 18782 2796 18788 2848
rect 18840 2836 18846 2848
rect 22830 2836 22836 2848
rect 18840 2808 22836 2836
rect 18840 2796 18846 2808
rect 22830 2796 22836 2808
rect 22888 2796 22894 2848
rect 28276 2836 28304 2876
rect 29917 2873 29929 2907
rect 29963 2904 29975 2907
rect 30282 2904 30288 2916
rect 29963 2876 30288 2904
rect 29963 2873 29975 2876
rect 29917 2867 29975 2873
rect 30282 2864 30288 2876
rect 30340 2864 30346 2916
rect 30374 2864 30380 2916
rect 30432 2904 30438 2916
rect 30852 2904 30880 2944
rect 32401 2941 32413 2975
rect 32447 2972 32459 2975
rect 32674 2972 32680 2984
rect 32447 2944 32680 2972
rect 32447 2941 32459 2944
rect 32401 2935 32459 2941
rect 32674 2932 32680 2944
rect 32732 2932 32738 2984
rect 32784 2981 32812 3012
rect 34330 3000 34336 3012
rect 34388 3000 34394 3052
rect 34606 3000 34612 3052
rect 34664 3040 34670 3052
rect 36096 3040 36124 3080
rect 36630 3068 36636 3080
rect 36688 3068 36694 3120
rect 34664 3012 36124 3040
rect 36449 3043 36507 3049
rect 34664 3000 34670 3012
rect 36449 3009 36461 3043
rect 36495 3040 36507 3043
rect 36722 3040 36728 3052
rect 36495 3012 36728 3040
rect 36495 3009 36507 3012
rect 36449 3003 36507 3009
rect 36722 3000 36728 3012
rect 36780 3000 36786 3052
rect 37936 3040 37964 3148
rect 38102 3136 38108 3188
rect 38160 3176 38166 3188
rect 39301 3179 39359 3185
rect 39301 3176 39313 3179
rect 38160 3148 39313 3176
rect 38160 3136 38166 3148
rect 39301 3145 39313 3148
rect 39347 3145 39359 3179
rect 39301 3139 39359 3145
rect 40662 3179 40720 3185
rect 40662 3145 40674 3179
rect 40708 3176 40720 3179
rect 41506 3176 41512 3188
rect 40708 3148 41512 3176
rect 40708 3145 40720 3148
rect 40662 3139 40720 3145
rect 38194 3040 38200 3052
rect 37936 3012 38056 3040
rect 38155 3012 38200 3040
rect 32769 2975 32827 2981
rect 32769 2941 32781 2975
rect 32815 2941 32827 2975
rect 32950 2972 32956 2984
rect 32911 2944 32956 2972
rect 32769 2935 32827 2941
rect 32950 2932 32956 2944
rect 33008 2932 33014 2984
rect 33781 2975 33839 2981
rect 33781 2941 33793 2975
rect 33827 2972 33839 2975
rect 35618 2972 35624 2984
rect 33827 2944 35624 2972
rect 33827 2941 33839 2944
rect 33781 2935 33839 2941
rect 35618 2932 35624 2944
rect 35676 2932 35682 2984
rect 35710 2932 35716 2984
rect 35768 2972 35774 2984
rect 37918 2972 37924 2984
rect 35768 2944 35813 2972
rect 36004 2944 36400 2972
rect 37879 2944 37924 2972
rect 35768 2932 35774 2944
rect 30432 2876 30880 2904
rect 30432 2864 30438 2876
rect 31386 2864 31392 2916
rect 31444 2904 31450 2916
rect 36004 2904 36032 2944
rect 31444 2876 36032 2904
rect 36081 2907 36139 2913
rect 31444 2864 31450 2876
rect 36081 2873 36093 2907
rect 36127 2904 36139 2907
rect 36262 2904 36268 2916
rect 36127 2876 36268 2904
rect 36127 2873 36139 2876
rect 36081 2867 36139 2873
rect 36262 2864 36268 2876
rect 36320 2864 36326 2916
rect 33042 2836 33048 2848
rect 28276 2808 33048 2836
rect 33042 2796 33048 2808
rect 33100 2796 33106 2848
rect 33873 2839 33931 2845
rect 33873 2805 33885 2839
rect 33919 2836 33931 2839
rect 35897 2839 35955 2845
rect 35897 2836 35909 2839
rect 33919 2808 35909 2836
rect 33919 2805 33931 2808
rect 33873 2799 33931 2805
rect 35897 2805 35909 2808
rect 35943 2805 35955 2839
rect 35897 2799 35955 2805
rect 35986 2796 35992 2848
rect 36044 2836 36050 2848
rect 36372 2836 36400 2944
rect 37918 2932 37924 2944
rect 37976 2932 37982 2984
rect 38028 2972 38056 3012
rect 38194 3000 38200 3012
rect 38252 3000 38258 3052
rect 39114 3040 39120 3052
rect 38396 3012 39120 3040
rect 38396 2972 38424 3012
rect 39114 3000 39120 3012
rect 39172 3000 39178 3052
rect 39316 3040 39344 3139
rect 41506 3136 41512 3148
rect 41564 3136 41570 3188
rect 44913 3179 44971 3185
rect 44913 3145 44925 3179
rect 44959 3176 44971 3179
rect 44959 3148 46796 3176
rect 44959 3145 44971 3148
rect 44913 3139 44971 3145
rect 40770 3108 40776 3120
rect 40731 3080 40776 3108
rect 40770 3068 40776 3080
rect 40828 3068 40834 3120
rect 46768 3108 46796 3148
rect 47026 3136 47032 3188
rect 47084 3176 47090 3188
rect 48574 3179 48632 3185
rect 48574 3176 48586 3179
rect 47084 3148 48586 3176
rect 47084 3136 47090 3148
rect 48574 3145 48586 3148
rect 48620 3176 48632 3179
rect 48620 3148 50384 3176
rect 48620 3145 48632 3148
rect 48574 3139 48632 3145
rect 48685 3111 48743 3117
rect 48685 3108 48697 3111
rect 46768 3080 48697 3108
rect 40865 3043 40923 3049
rect 40865 3040 40877 3043
rect 39316 3012 40877 3040
rect 40865 3009 40877 3012
rect 40911 3009 40923 3043
rect 40865 3003 40923 3009
rect 41233 3043 41291 3049
rect 41233 3009 41245 3043
rect 41279 3040 41291 3043
rect 41279 3012 46152 3040
rect 41279 3009 41291 3012
rect 41233 3003 41291 3009
rect 38028 2944 38424 2972
rect 38470 2932 38476 2984
rect 38528 2972 38534 2984
rect 40880 2972 40908 3003
rect 41322 2972 41328 2984
rect 38528 2944 40632 2972
rect 40880 2944 41328 2972
rect 38528 2932 38534 2944
rect 40494 2904 40500 2916
rect 40455 2876 40500 2904
rect 40494 2864 40500 2876
rect 40552 2864 40558 2916
rect 40604 2904 40632 2944
rect 41322 2932 41328 2944
rect 41380 2932 41386 2984
rect 42058 2972 42064 2984
rect 42019 2944 42064 2972
rect 42058 2932 42064 2944
rect 42116 2932 42122 2984
rect 44821 2975 44879 2981
rect 44821 2941 44833 2975
rect 44867 2972 44879 2975
rect 45186 2972 45192 2984
rect 44867 2944 45192 2972
rect 44867 2941 44879 2944
rect 44821 2935 44879 2941
rect 45186 2932 45192 2944
rect 45244 2932 45250 2984
rect 46124 2981 46152 3012
rect 46768 2981 46796 3080
rect 48685 3077 48697 3080
rect 48731 3077 48743 3111
rect 50356 3108 50384 3148
rect 51258 3136 51264 3188
rect 51316 3176 51322 3188
rect 52454 3176 52460 3188
rect 51316 3148 52460 3176
rect 51316 3136 51322 3148
rect 52454 3136 52460 3148
rect 52512 3136 52518 3188
rect 53466 3176 53472 3188
rect 53427 3148 53472 3176
rect 53466 3136 53472 3148
rect 53524 3136 53530 3188
rect 53558 3136 53564 3188
rect 53616 3176 53622 3188
rect 58483 3179 58541 3185
rect 58483 3176 58495 3179
rect 53616 3148 58495 3176
rect 53616 3136 53622 3148
rect 58483 3145 58495 3148
rect 58529 3145 58541 3179
rect 58483 3139 58541 3145
rect 57974 3108 57980 3120
rect 50356 3080 57980 3108
rect 48685 3071 48743 3077
rect 57974 3068 57980 3080
rect 58032 3068 58038 3120
rect 58621 3111 58679 3117
rect 58621 3077 58633 3111
rect 58667 3108 58679 3111
rect 61930 3108 61936 3120
rect 58667 3080 61936 3108
rect 58667 3077 58679 3080
rect 58621 3071 58679 3077
rect 61930 3068 61936 3080
rect 61988 3068 61994 3120
rect 48777 3043 48835 3049
rect 48777 3040 48789 3043
rect 47320 3012 48789 3040
rect 46109 2975 46167 2981
rect 46109 2941 46121 2975
rect 46155 2941 46167 2975
rect 46109 2935 46167 2941
rect 46753 2975 46811 2981
rect 46753 2941 46765 2975
rect 46799 2941 46811 2975
rect 47026 2972 47032 2984
rect 46987 2944 47032 2972
rect 46753 2935 46811 2941
rect 42153 2907 42211 2913
rect 42153 2904 42165 2907
rect 40604 2876 42165 2904
rect 42153 2873 42165 2876
rect 42199 2873 42211 2907
rect 44634 2904 44640 2916
rect 44595 2876 44640 2904
rect 42153 2867 42211 2873
rect 44634 2864 44640 2876
rect 44692 2864 44698 2916
rect 46124 2904 46152 2935
rect 47026 2932 47032 2944
rect 47084 2932 47090 2984
rect 46124 2876 46796 2904
rect 43346 2836 43352 2848
rect 36044 2808 36089 2836
rect 36372 2808 43352 2836
rect 36044 2796 36050 2808
rect 43346 2796 43352 2808
rect 43404 2796 43410 2848
rect 44082 2796 44088 2848
rect 44140 2836 44146 2848
rect 46201 2839 46259 2845
rect 46201 2836 46213 2839
rect 44140 2808 46213 2836
rect 44140 2796 44146 2808
rect 46201 2805 46213 2808
rect 46247 2805 46259 2839
rect 46768 2836 46796 2876
rect 47320 2836 47348 3012
rect 48777 3009 48789 3012
rect 48823 3009 48835 3043
rect 48777 3003 48835 3009
rect 52178 3000 52184 3052
rect 52236 3040 52242 3052
rect 53929 3043 53987 3049
rect 53929 3040 53941 3043
rect 52236 3012 53941 3040
rect 52236 3000 52242 3012
rect 53929 3009 53941 3012
rect 53975 3009 53987 3043
rect 53929 3003 53987 3009
rect 55398 3000 55404 3052
rect 55456 3040 55462 3052
rect 55861 3043 55919 3049
rect 55861 3040 55873 3043
rect 55456 3012 55873 3040
rect 55456 3000 55462 3012
rect 55861 3009 55873 3012
rect 55907 3009 55919 3043
rect 58710 3040 58716 3052
rect 58671 3012 58716 3040
rect 55861 3003 55919 3009
rect 58710 3000 58716 3012
rect 58768 3000 58774 3052
rect 47489 2975 47547 2981
rect 47489 2941 47501 2975
rect 47535 2941 47547 2975
rect 47489 2935 47547 2941
rect 47504 2904 47532 2935
rect 47578 2932 47584 2984
rect 47636 2972 47642 2984
rect 49786 2972 49792 2984
rect 47636 2944 49792 2972
rect 47636 2932 47642 2944
rect 49786 2932 49792 2944
rect 49844 2932 49850 2984
rect 49970 2972 49976 2984
rect 49931 2944 49976 2972
rect 49970 2932 49976 2944
rect 50028 2932 50034 2984
rect 52273 2975 52331 2981
rect 52273 2941 52285 2975
rect 52319 2972 52331 2975
rect 53742 2972 53748 2984
rect 52319 2944 53748 2972
rect 52319 2941 52331 2944
rect 52273 2935 52331 2941
rect 53742 2932 53748 2944
rect 53800 2932 53806 2984
rect 54018 2972 54024 2984
rect 53979 2944 54024 2972
rect 54018 2932 54024 2944
rect 54076 2932 54082 2984
rect 54386 2972 54392 2984
rect 54347 2944 54392 2972
rect 54386 2932 54392 2944
rect 54444 2932 54450 2984
rect 54570 2972 54576 2984
rect 54531 2944 54576 2972
rect 54570 2932 54576 2944
rect 54628 2932 54634 2984
rect 54662 2932 54668 2984
rect 54720 2972 54726 2984
rect 55582 2972 55588 2984
rect 54720 2944 55444 2972
rect 55543 2944 55588 2972
rect 54720 2932 54726 2944
rect 55416 2913 55444 2944
rect 55582 2932 55588 2944
rect 55640 2932 55646 2984
rect 56686 2932 56692 2984
rect 56744 2972 56750 2984
rect 60093 2975 60151 2981
rect 60093 2972 60105 2975
rect 56744 2944 60105 2972
rect 56744 2932 56750 2944
rect 60093 2941 60105 2944
rect 60139 2941 60151 2975
rect 60093 2935 60151 2941
rect 48409 2907 48467 2913
rect 48409 2904 48421 2907
rect 47504 2876 48421 2904
rect 48409 2873 48421 2876
rect 48455 2904 48467 2907
rect 55401 2907 55459 2913
rect 48455 2876 55352 2904
rect 48455 2873 48467 2876
rect 48409 2867 48467 2873
rect 46768 2808 47348 2836
rect 46201 2799 46259 2805
rect 48498 2796 48504 2848
rect 48556 2836 48562 2848
rect 49053 2839 49111 2845
rect 49053 2836 49065 2839
rect 48556 2808 49065 2836
rect 48556 2796 48562 2808
rect 49053 2805 49065 2808
rect 49099 2805 49111 2839
rect 49053 2799 49111 2805
rect 49786 2796 49792 2848
rect 49844 2836 49850 2848
rect 50157 2839 50215 2845
rect 50157 2836 50169 2839
rect 49844 2808 50169 2836
rect 49844 2796 49850 2808
rect 50157 2805 50169 2808
rect 50203 2836 50215 2839
rect 54662 2836 54668 2848
rect 50203 2808 54668 2836
rect 50203 2805 50215 2808
rect 50157 2799 50215 2805
rect 54662 2796 54668 2808
rect 54720 2796 54726 2848
rect 55324 2836 55352 2876
rect 55401 2873 55413 2907
rect 55447 2904 55459 2907
rect 56778 2904 56784 2916
rect 55447 2876 56784 2904
rect 55447 2873 55459 2876
rect 55401 2867 55459 2873
rect 56778 2864 56784 2876
rect 56836 2864 56842 2916
rect 58345 2907 58403 2913
rect 58345 2873 58357 2907
rect 58391 2904 58403 2907
rect 58391 2876 59216 2904
rect 58391 2873 58403 2876
rect 58345 2867 58403 2873
rect 58989 2839 59047 2845
rect 58989 2836 59001 2839
rect 55324 2808 59001 2836
rect 58989 2805 59001 2808
rect 59035 2805 59047 2839
rect 59188 2836 59216 2876
rect 59262 2864 59268 2916
rect 59320 2904 59326 2916
rect 59909 2907 59967 2913
rect 59909 2904 59921 2907
rect 59320 2876 59921 2904
rect 59320 2864 59326 2876
rect 59909 2873 59921 2876
rect 59955 2873 59967 2907
rect 59909 2867 59967 2873
rect 60185 2839 60243 2845
rect 60185 2836 60197 2839
rect 59188 2808 60197 2836
rect 58989 2799 59047 2805
rect 60185 2805 60197 2808
rect 60231 2805 60243 2839
rect 60185 2799 60243 2805
rect 60642 2796 60648 2848
rect 60700 2836 60706 2848
rect 62758 2836 62764 2848
rect 60700 2808 62764 2836
rect 60700 2796 60706 2808
rect 62758 2796 62764 2808
rect 62816 2796 62822 2848
rect 1104 2746 62192 2768
rect 1104 2694 21344 2746
rect 21396 2694 21408 2746
rect 21460 2694 21472 2746
rect 21524 2694 21536 2746
rect 21588 2694 41707 2746
rect 41759 2694 41771 2746
rect 41823 2694 41835 2746
rect 41887 2694 41899 2746
rect 41951 2694 62192 2746
rect 1104 2672 62192 2694
rect 22094 2632 22100 2644
rect 2792 2604 22100 2632
rect 2038 2456 2044 2508
rect 2096 2496 2102 2508
rect 2792 2505 2820 2604
rect 22094 2592 22100 2604
rect 22152 2592 22158 2644
rect 30006 2592 30012 2644
rect 30064 2632 30070 2644
rect 35529 2635 35587 2641
rect 35529 2632 35541 2635
rect 30064 2604 35541 2632
rect 30064 2592 30070 2604
rect 5997 2567 6055 2573
rect 5997 2533 6009 2567
rect 6043 2564 6055 2567
rect 6822 2564 6828 2576
rect 6043 2536 6828 2564
rect 6043 2533 6055 2536
rect 5997 2527 6055 2533
rect 6822 2524 6828 2536
rect 6880 2524 6886 2576
rect 8573 2567 8631 2573
rect 8573 2533 8585 2567
rect 8619 2564 8631 2567
rect 8662 2564 8668 2576
rect 8619 2536 8668 2564
rect 8619 2533 8631 2536
rect 8573 2527 8631 2533
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 20806 2524 20812 2576
rect 20864 2564 20870 2576
rect 21361 2567 21419 2573
rect 21361 2564 21373 2567
rect 20864 2536 21373 2564
rect 20864 2524 20870 2536
rect 21361 2533 21373 2536
rect 21407 2533 21419 2567
rect 21361 2527 21419 2533
rect 25961 2567 26019 2573
rect 25961 2533 25973 2567
rect 26007 2564 26019 2567
rect 26050 2564 26056 2576
rect 26007 2536 26056 2564
rect 26007 2533 26019 2536
rect 25961 2527 26019 2533
rect 26050 2524 26056 2536
rect 26108 2524 26114 2576
rect 26160 2536 27660 2564
rect 2409 2499 2467 2505
rect 2409 2496 2421 2499
rect 2096 2468 2421 2496
rect 2096 2456 2102 2468
rect 2409 2465 2421 2468
rect 2455 2465 2467 2499
rect 2409 2459 2467 2465
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2465 2835 2499
rect 2958 2496 2964 2508
rect 2919 2468 2964 2496
rect 2777 2459 2835 2465
rect 2958 2456 2964 2468
rect 3016 2456 3022 2508
rect 4617 2499 4675 2505
rect 4617 2465 4629 2499
rect 4663 2496 4675 2499
rect 5534 2496 5540 2508
rect 4663 2468 5540 2496
rect 4663 2465 4675 2468
rect 4617 2459 4675 2465
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 5902 2456 5908 2508
rect 5960 2496 5966 2508
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 5960 2468 7205 2496
rect 5960 2456 5966 2468
rect 7193 2465 7205 2468
rect 7239 2465 7251 2499
rect 7193 2459 7251 2465
rect 12342 2456 12348 2508
rect 12400 2496 12406 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12400 2468 12633 2496
rect 12400 2456 12406 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12894 2496 12900 2508
rect 12855 2468 12900 2496
rect 12621 2459 12679 2465
rect 12894 2456 12900 2468
rect 12952 2456 12958 2508
rect 16025 2499 16083 2505
rect 16025 2465 16037 2499
rect 16071 2496 16083 2499
rect 17310 2496 17316 2508
rect 16071 2468 17316 2496
rect 16071 2465 16083 2468
rect 16025 2459 16083 2465
rect 17310 2456 17316 2468
rect 17368 2456 17374 2508
rect 17586 2456 17592 2508
rect 17644 2496 17650 2508
rect 18601 2499 18659 2505
rect 18601 2496 18613 2499
rect 17644 2468 18613 2496
rect 17644 2456 17650 2468
rect 18601 2465 18613 2468
rect 18647 2465 18659 2499
rect 18601 2459 18659 2465
rect 21082 2456 21088 2508
rect 21140 2496 21146 2508
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 21140 2468 21189 2496
rect 21140 2456 21146 2468
rect 21177 2465 21189 2468
rect 21223 2465 21235 2499
rect 21177 2459 21235 2465
rect 21453 2499 21511 2505
rect 21453 2465 21465 2499
rect 21499 2465 21511 2499
rect 21453 2459 21511 2465
rect 4338 2428 4344 2440
rect 4251 2400 4344 2428
rect 4338 2388 4344 2400
rect 4396 2428 4402 2440
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 4396 2400 6929 2428
rect 4396 2388 4402 2400
rect 6917 2397 6929 2400
rect 6963 2428 6975 2431
rect 12360 2428 12388 2456
rect 6963 2400 12388 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 14001 2431 14059 2437
rect 14001 2428 14013 2431
rect 12860 2400 14013 2428
rect 12860 2388 12866 2400
rect 14001 2397 14013 2400
rect 14047 2397 14059 2431
rect 14001 2391 14059 2397
rect 15749 2431 15807 2437
rect 15749 2397 15761 2431
rect 15795 2428 15807 2431
rect 16390 2428 16396 2440
rect 15795 2400 16396 2428
rect 15795 2397 15807 2400
rect 15749 2391 15807 2397
rect 16390 2388 16396 2400
rect 16448 2388 16454 2440
rect 16666 2388 16672 2440
rect 16724 2428 16730 2440
rect 17129 2431 17187 2437
rect 17129 2428 17141 2431
rect 16724 2400 17141 2428
rect 16724 2388 16730 2400
rect 17129 2397 17141 2400
rect 17175 2397 17187 2431
rect 18322 2428 18328 2440
rect 18283 2400 18328 2428
rect 17129 2391 17187 2397
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 19702 2428 19708 2440
rect 19663 2400 19708 2428
rect 19702 2388 19708 2400
rect 19760 2388 19766 2440
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 21468 2428 21496 2459
rect 22830 2456 22836 2508
rect 22888 2496 22894 2508
rect 22925 2499 22983 2505
rect 22925 2496 22937 2499
rect 22888 2468 22937 2496
rect 22888 2456 22894 2468
rect 22925 2465 22937 2468
rect 22971 2465 22983 2499
rect 22925 2459 22983 2465
rect 23017 2499 23075 2505
rect 23017 2465 23029 2499
rect 23063 2496 23075 2499
rect 26160 2496 26188 2536
rect 26878 2496 26884 2508
rect 23063 2468 26188 2496
rect 26839 2468 26884 2496
rect 23063 2465 23075 2468
rect 23017 2459 23075 2465
rect 26878 2456 26884 2468
rect 26936 2456 26942 2508
rect 27632 2505 27660 2536
rect 31018 2524 31024 2576
rect 31076 2564 31082 2576
rect 32582 2564 32588 2576
rect 31076 2536 32588 2564
rect 31076 2524 31082 2536
rect 32582 2524 32588 2536
rect 32640 2524 32646 2576
rect 27617 2499 27675 2505
rect 27617 2465 27629 2499
rect 27663 2465 27675 2499
rect 27617 2459 27675 2465
rect 28077 2499 28135 2505
rect 28077 2465 28089 2499
rect 28123 2496 28135 2499
rect 28258 2496 28264 2508
rect 28123 2468 28264 2496
rect 28123 2465 28135 2468
rect 28077 2459 28135 2465
rect 28258 2456 28264 2468
rect 28316 2456 28322 2508
rect 30282 2496 30288 2508
rect 30243 2468 30288 2496
rect 30282 2456 30288 2468
rect 30340 2456 30346 2508
rect 32692 2505 32720 2604
rect 35529 2601 35541 2604
rect 35575 2601 35587 2635
rect 35529 2595 35587 2601
rect 41506 2592 41512 2644
rect 41564 2632 41570 2644
rect 41785 2635 41843 2641
rect 41785 2632 41797 2635
rect 41564 2604 41797 2632
rect 41564 2592 41570 2604
rect 41785 2601 41797 2604
rect 41831 2601 41843 2635
rect 41785 2595 41843 2601
rect 44634 2592 44640 2644
rect 44692 2632 44698 2644
rect 45097 2635 45155 2641
rect 45097 2632 45109 2635
rect 44692 2604 45109 2632
rect 44692 2592 44698 2604
rect 45097 2601 45109 2604
rect 45143 2601 45155 2635
rect 45097 2595 45155 2601
rect 45186 2592 45192 2644
rect 45244 2632 45250 2644
rect 47581 2635 47639 2641
rect 47581 2632 47593 2635
rect 45244 2604 47593 2632
rect 45244 2592 45250 2604
rect 47581 2601 47593 2604
rect 47627 2601 47639 2635
rect 47581 2595 47639 2601
rect 48590 2592 48596 2644
rect 48648 2632 48654 2644
rect 48685 2635 48743 2641
rect 48685 2632 48697 2635
rect 48648 2604 48697 2632
rect 48648 2592 48654 2604
rect 48685 2601 48697 2604
rect 48731 2601 48743 2635
rect 48685 2595 48743 2601
rect 57974 2592 57980 2644
rect 58032 2632 58038 2644
rect 58897 2635 58955 2641
rect 58897 2632 58909 2635
rect 58032 2604 58909 2632
rect 58032 2592 58038 2604
rect 58897 2601 58909 2604
rect 58943 2601 58955 2635
rect 58897 2595 58955 2601
rect 33962 2564 33968 2576
rect 33923 2536 33968 2564
rect 33962 2524 33968 2536
rect 34020 2524 34026 2576
rect 38102 2564 38108 2576
rect 34164 2536 38108 2564
rect 34164 2505 34192 2536
rect 38102 2524 38108 2536
rect 38160 2524 38166 2576
rect 40221 2567 40279 2573
rect 40221 2533 40233 2567
rect 40267 2564 40279 2567
rect 40770 2564 40776 2576
rect 40267 2536 40776 2564
rect 40267 2533 40279 2536
rect 40221 2527 40279 2533
rect 40770 2524 40776 2536
rect 40828 2524 40834 2576
rect 56781 2567 56839 2573
rect 56781 2533 56793 2567
rect 56827 2564 56839 2567
rect 58434 2564 58440 2576
rect 56827 2536 58440 2564
rect 56827 2533 56839 2536
rect 56781 2527 56839 2533
rect 58434 2524 58440 2536
rect 58492 2524 58498 2576
rect 32677 2499 32735 2505
rect 32677 2465 32689 2499
rect 32723 2465 32735 2499
rect 32677 2459 32735 2465
rect 34149 2499 34207 2505
rect 34149 2465 34161 2499
rect 34195 2465 34207 2499
rect 34149 2459 34207 2465
rect 35713 2499 35771 2505
rect 35713 2465 35725 2499
rect 35759 2465 35771 2499
rect 35894 2496 35900 2508
rect 35855 2468 35900 2496
rect 35713 2459 35771 2465
rect 24302 2428 24308 2440
rect 20772 2400 21496 2428
rect 24215 2400 24308 2428
rect 20772 2388 20778 2400
rect 24302 2388 24308 2400
rect 24360 2388 24366 2440
rect 24581 2431 24639 2437
rect 24581 2397 24593 2431
rect 24627 2428 24639 2431
rect 30009 2431 30067 2437
rect 30009 2428 30021 2431
rect 24627 2400 27200 2428
rect 24627 2397 24639 2400
rect 24581 2391 24639 2397
rect 17954 2252 17960 2304
rect 18012 2292 18018 2304
rect 21637 2295 21695 2301
rect 21637 2292 21649 2295
rect 18012 2264 21649 2292
rect 18012 2252 18018 2264
rect 21637 2261 21649 2264
rect 21683 2261 21695 2295
rect 21637 2255 21695 2261
rect 21726 2252 21732 2304
rect 21784 2292 21790 2304
rect 24320 2292 24348 2388
rect 27172 2369 27200 2400
rect 27264 2400 30021 2428
rect 27157 2363 27215 2369
rect 27157 2329 27169 2363
rect 27203 2329 27215 2363
rect 27157 2323 27215 2329
rect 24946 2292 24952 2304
rect 21784 2264 24952 2292
rect 21784 2252 21790 2264
rect 24946 2252 24952 2264
rect 25004 2292 25010 2304
rect 27264 2292 27292 2400
rect 30009 2397 30021 2400
rect 30055 2397 30067 2431
rect 30009 2391 30067 2397
rect 31110 2388 31116 2440
rect 31168 2428 31174 2440
rect 32585 2431 32643 2437
rect 32585 2428 32597 2431
rect 31168 2400 32597 2428
rect 31168 2388 31174 2400
rect 32585 2397 32597 2400
rect 32631 2428 32643 2431
rect 32766 2428 32772 2440
rect 32631 2400 32772 2428
rect 32631 2397 32643 2400
rect 32585 2391 32643 2397
rect 32766 2388 32772 2400
rect 32824 2388 32830 2440
rect 34517 2431 34575 2437
rect 34517 2397 34529 2431
rect 34563 2428 34575 2431
rect 34606 2428 34612 2440
rect 34563 2400 34612 2428
rect 34563 2397 34575 2400
rect 34517 2391 34575 2397
rect 34606 2388 34612 2400
rect 34664 2388 34670 2440
rect 35728 2428 35756 2459
rect 35894 2456 35900 2468
rect 35952 2456 35958 2508
rect 36262 2496 36268 2508
rect 36223 2468 36268 2496
rect 36262 2456 36268 2468
rect 36320 2456 36326 2508
rect 37918 2456 37924 2508
rect 37976 2496 37982 2508
rect 38565 2499 38623 2505
rect 38565 2496 38577 2499
rect 37976 2468 38577 2496
rect 37976 2456 37982 2468
rect 38565 2465 38577 2468
rect 38611 2465 38623 2499
rect 38565 2459 38623 2465
rect 38654 2456 38660 2508
rect 38712 2496 38718 2508
rect 38841 2499 38899 2505
rect 38841 2496 38853 2499
rect 38712 2468 38853 2496
rect 38712 2456 38718 2468
rect 38841 2465 38853 2468
rect 38887 2465 38899 2499
rect 38841 2459 38899 2465
rect 41046 2456 41052 2508
rect 41104 2496 41110 2508
rect 41141 2499 41199 2505
rect 41141 2496 41153 2499
rect 41104 2468 41153 2496
rect 41104 2456 41110 2468
rect 41141 2465 41153 2468
rect 41187 2465 41199 2499
rect 41141 2459 41199 2465
rect 41322 2456 41328 2508
rect 41380 2496 41386 2508
rect 42705 2499 42763 2505
rect 42705 2496 42717 2499
rect 41380 2468 42717 2496
rect 41380 2456 41386 2468
rect 42705 2465 42717 2468
rect 42751 2465 42763 2499
rect 42705 2459 42763 2465
rect 44453 2499 44511 2505
rect 44453 2465 44465 2499
rect 44499 2496 44511 2499
rect 44542 2496 44548 2508
rect 44499 2468 44548 2496
rect 44499 2465 44511 2468
rect 44453 2459 44511 2465
rect 44542 2456 44548 2468
rect 44600 2456 44606 2508
rect 46937 2499 46995 2505
rect 46937 2465 46949 2499
rect 46983 2496 46995 2499
rect 48038 2496 48044 2508
rect 46983 2468 48044 2496
rect 46983 2465 46995 2468
rect 46937 2459 46995 2465
rect 48038 2456 48044 2468
rect 48096 2456 48102 2508
rect 48498 2496 48504 2508
rect 48459 2468 48504 2496
rect 48498 2456 48504 2468
rect 48556 2456 48562 2508
rect 53745 2499 53803 2505
rect 53745 2465 53757 2499
rect 53791 2496 53803 2499
rect 54938 2496 54944 2508
rect 53791 2468 54944 2496
rect 53791 2465 53803 2468
rect 53745 2459 53803 2465
rect 54938 2456 54944 2468
rect 54996 2456 55002 2508
rect 56965 2499 57023 2505
rect 56965 2465 56977 2499
rect 57011 2465 57023 2499
rect 56965 2459 57023 2465
rect 57333 2499 57391 2505
rect 57333 2465 57345 2499
rect 57379 2496 57391 2499
rect 58253 2499 58311 2505
rect 58253 2496 58265 2499
rect 57379 2468 58265 2496
rect 57379 2465 57391 2468
rect 57333 2459 57391 2465
rect 58253 2465 58265 2468
rect 58299 2465 58311 2499
rect 58253 2459 58311 2465
rect 59817 2499 59875 2505
rect 59817 2465 59829 2499
rect 59863 2496 59875 2499
rect 60182 2496 60188 2508
rect 59863 2468 60188 2496
rect 59863 2465 59875 2468
rect 59817 2459 59875 2465
rect 36078 2428 36084 2440
rect 35728 2400 36084 2428
rect 36078 2388 36084 2400
rect 36136 2388 36142 2440
rect 40218 2388 40224 2440
rect 40276 2428 40282 2440
rect 41509 2431 41567 2437
rect 41509 2428 41521 2431
rect 40276 2400 41521 2428
rect 40276 2388 40282 2400
rect 41509 2397 41521 2400
rect 41555 2397 41567 2431
rect 41509 2391 41567 2397
rect 43714 2388 43720 2440
rect 43772 2428 43778 2440
rect 44821 2431 44879 2437
rect 44821 2428 44833 2431
rect 43772 2400 44833 2428
rect 43772 2388 43778 2400
rect 44821 2397 44833 2400
rect 44867 2397 44879 2431
rect 44821 2391 44879 2397
rect 47118 2388 47124 2440
rect 47176 2428 47182 2440
rect 47305 2431 47363 2437
rect 47305 2428 47317 2431
rect 47176 2400 47317 2428
rect 47176 2388 47182 2400
rect 47305 2397 47317 2400
rect 47351 2397 47363 2431
rect 47305 2391 47363 2397
rect 49786 2388 49792 2440
rect 49844 2428 49850 2440
rect 54113 2431 54171 2437
rect 54113 2428 54125 2431
rect 49844 2400 54125 2428
rect 49844 2388 49850 2400
rect 54113 2397 54125 2400
rect 54159 2397 54171 2431
rect 56980 2428 57008 2459
rect 60182 2456 60188 2468
rect 60240 2456 60246 2508
rect 57606 2428 57612 2440
rect 56980 2400 57612 2428
rect 54113 2391 54171 2397
rect 57606 2388 57612 2400
rect 57664 2388 57670 2440
rect 58621 2431 58679 2437
rect 58621 2397 58633 2431
rect 58667 2428 58679 2431
rect 59909 2431 59967 2437
rect 59909 2428 59921 2431
rect 58667 2400 59921 2428
rect 58667 2397 58679 2400
rect 58621 2391 58679 2397
rect 59909 2397 59921 2400
rect 59955 2397 59967 2431
rect 59909 2391 59967 2397
rect 41306 2363 41364 2369
rect 41306 2329 41318 2363
rect 41352 2360 41364 2363
rect 41966 2360 41972 2372
rect 41352 2332 41972 2360
rect 41352 2329 41364 2332
rect 41306 2323 41364 2329
rect 41966 2320 41972 2332
rect 42024 2320 42030 2372
rect 44618 2363 44676 2369
rect 44618 2329 44630 2363
rect 44664 2360 44676 2363
rect 45462 2360 45468 2372
rect 44664 2332 45468 2360
rect 44664 2329 44676 2332
rect 44618 2323 44676 2329
rect 45462 2320 45468 2332
rect 45520 2320 45526 2372
rect 46290 2320 46296 2372
rect 46348 2360 46354 2372
rect 47213 2363 47271 2369
rect 47213 2360 47225 2363
rect 46348 2332 47225 2360
rect 46348 2320 46354 2332
rect 47213 2329 47225 2332
rect 47259 2329 47271 2363
rect 47213 2323 47271 2329
rect 53910 2363 53968 2369
rect 53910 2329 53922 2363
rect 53956 2360 53968 2363
rect 54389 2363 54447 2369
rect 53956 2332 54156 2360
rect 53956 2329 53968 2332
rect 53910 2323 53968 2329
rect 54128 2304 54156 2332
rect 54389 2329 54401 2363
rect 54435 2360 54447 2363
rect 58391 2363 58449 2369
rect 58391 2360 58403 2363
rect 54435 2332 58403 2360
rect 54435 2329 54447 2332
rect 54389 2323 54447 2329
rect 58391 2329 58403 2332
rect 58437 2329 58449 2363
rect 58391 2323 58449 2329
rect 58529 2363 58587 2369
rect 58529 2329 58541 2363
rect 58575 2360 58587 2363
rect 60642 2360 60648 2372
rect 58575 2332 60648 2360
rect 58575 2329 58587 2332
rect 58529 2323 58587 2329
rect 60642 2320 60648 2332
rect 60700 2320 60706 2372
rect 25004 2264 27292 2292
rect 25004 2252 25010 2264
rect 29730 2252 29736 2304
rect 29788 2292 29794 2304
rect 31389 2295 31447 2301
rect 31389 2292 31401 2295
rect 29788 2264 31401 2292
rect 29788 2252 29794 2264
rect 31389 2261 31401 2264
rect 31435 2261 31447 2295
rect 32858 2292 32864 2304
rect 32819 2264 32864 2292
rect 31389 2255 31447 2261
rect 32858 2252 32864 2264
rect 32916 2252 32922 2304
rect 39482 2252 39488 2304
rect 39540 2292 39546 2304
rect 41417 2295 41475 2301
rect 41417 2292 41429 2295
rect 39540 2264 41429 2292
rect 39540 2252 39546 2264
rect 41417 2261 41429 2264
rect 41463 2261 41475 2295
rect 42794 2292 42800 2304
rect 42755 2264 42800 2292
rect 41417 2255 41475 2261
rect 42794 2252 42800 2264
rect 42852 2252 42858 2304
rect 42886 2252 42892 2304
rect 42944 2292 42950 2304
rect 44729 2295 44787 2301
rect 44729 2292 44741 2295
rect 42944 2264 44741 2292
rect 42944 2252 42950 2264
rect 44729 2261 44741 2264
rect 44775 2261 44787 2295
rect 44729 2255 44787 2261
rect 47102 2295 47160 2301
rect 47102 2261 47114 2295
rect 47148 2292 47160 2295
rect 48866 2292 48872 2304
rect 47148 2264 48872 2292
rect 47148 2261 47160 2264
rect 47102 2255 47160 2261
rect 48866 2252 48872 2264
rect 48924 2252 48930 2304
rect 52362 2252 52368 2304
rect 52420 2292 52426 2304
rect 54021 2295 54079 2301
rect 54021 2292 54033 2295
rect 52420 2264 54033 2292
rect 52420 2252 52426 2264
rect 54021 2261 54033 2264
rect 54067 2261 54079 2295
rect 54021 2255 54079 2261
rect 54110 2252 54116 2304
rect 54168 2252 54174 2304
rect 1104 2202 62192 2224
rect 1104 2150 11163 2202
rect 11215 2150 11227 2202
rect 11279 2150 11291 2202
rect 11343 2150 11355 2202
rect 11407 2150 31526 2202
rect 31578 2150 31590 2202
rect 31642 2150 31654 2202
rect 31706 2150 31718 2202
rect 31770 2150 51888 2202
rect 51940 2150 51952 2202
rect 52004 2150 52016 2202
rect 52068 2150 52080 2202
rect 52132 2150 62192 2202
rect 1104 2128 62192 2150
rect 16390 2048 16396 2100
rect 16448 2088 16454 2100
rect 18322 2088 18328 2100
rect 16448 2060 18328 2088
rect 16448 2048 16454 2060
rect 18322 2048 18328 2060
rect 18380 2088 18386 2100
rect 21726 2088 21732 2100
rect 18380 2060 21732 2088
rect 18380 2048 18386 2060
rect 21726 2048 21732 2060
rect 21784 2048 21790 2100
rect 22094 2048 22100 2100
rect 22152 2088 22158 2100
rect 31018 2088 31024 2100
rect 22152 2060 31024 2088
rect 22152 2048 22158 2060
rect 31018 2048 31024 2060
rect 31076 2048 31082 2100
rect 32582 2048 32588 2100
rect 32640 2088 32646 2100
rect 40494 2088 40500 2100
rect 32640 2060 40500 2088
rect 32640 2048 32646 2060
rect 40494 2048 40500 2060
rect 40552 2048 40558 2100
rect 14458 1980 14464 2032
rect 14516 2020 14522 2032
rect 16850 2020 16856 2032
rect 14516 1992 16856 2020
rect 14516 1980 14522 1992
rect 16850 1980 16856 1992
rect 16908 1980 16914 2032
rect 36262 1980 36268 2032
rect 36320 2020 36326 2032
rect 37642 2020 37648 2032
rect 36320 1992 37648 2020
rect 36320 1980 36326 1992
rect 37642 1980 37648 1992
rect 37700 1980 37706 2032
rect 42794 2020 42800 2032
rect 38580 1992 42800 2020
rect 12710 1912 12716 1964
rect 12768 1952 12774 1964
rect 13354 1952 13360 1964
rect 12768 1924 13360 1952
rect 12768 1912 12774 1924
rect 13354 1912 13360 1924
rect 13412 1952 13418 1964
rect 18966 1952 18972 1964
rect 13412 1924 18972 1952
rect 13412 1912 13418 1924
rect 18966 1912 18972 1924
rect 19024 1912 19030 1964
rect 36354 1912 36360 1964
rect 36412 1952 36418 1964
rect 38580 1952 38608 1992
rect 42794 1980 42800 1992
rect 42852 1980 42858 2032
rect 36412 1924 38608 1952
rect 36412 1912 36418 1924
rect 32766 1844 32772 1896
rect 32824 1884 32830 1896
rect 34790 1884 34796 1896
rect 32824 1856 34796 1884
rect 32824 1844 32830 1856
rect 34790 1844 34796 1856
rect 34848 1884 34854 1896
rect 38470 1884 38476 1896
rect 34848 1856 38476 1884
rect 34848 1844 34854 1856
rect 38470 1844 38476 1856
rect 38528 1844 38534 1896
rect 36078 1776 36084 1828
rect 36136 1816 36142 1828
rect 36722 1816 36728 1828
rect 36136 1788 36728 1816
rect 36136 1776 36142 1788
rect 36722 1776 36728 1788
rect 36780 1776 36786 1828
rect 3418 1300 3424 1352
rect 3476 1340 3482 1352
rect 27154 1340 27160 1352
rect 3476 1312 27160 1340
rect 3476 1300 3482 1312
rect 27154 1300 27160 1312
rect 27212 1300 27218 1352
<< via1 >>
rect 11163 17382 11215 17434
rect 11227 17382 11279 17434
rect 11291 17382 11343 17434
rect 11355 17382 11407 17434
rect 31526 17382 31578 17434
rect 31590 17382 31642 17434
rect 31654 17382 31706 17434
rect 31718 17382 31770 17434
rect 51888 17382 51940 17434
rect 51952 17382 52004 17434
rect 52016 17382 52068 17434
rect 52080 17382 52132 17434
rect 14372 17323 14424 17332
rect 14372 17289 14381 17323
rect 14381 17289 14415 17323
rect 14415 17289 14424 17323
rect 14372 17280 14424 17289
rect 16212 17280 16264 17332
rect 20076 17280 20128 17332
rect 25412 17280 25464 17332
rect 27712 17280 27764 17332
rect 40500 17280 40552 17332
rect 41144 17280 41196 17332
rect 45008 17280 45060 17332
rect 11704 17144 11756 17196
rect 16672 17144 16724 17196
rect 13084 17119 13136 17128
rect 13084 17085 13093 17119
rect 13093 17085 13127 17119
rect 13127 17085 13136 17119
rect 13084 17076 13136 17085
rect 17960 17076 18012 17128
rect 18420 17076 18472 17128
rect 18604 17119 18656 17128
rect 18604 17085 18613 17119
rect 18613 17085 18647 17119
rect 18647 17085 18656 17119
rect 18604 17076 18656 17085
rect 25872 17144 25924 17196
rect 24032 17119 24084 17128
rect 24032 17085 24041 17119
rect 24041 17085 24075 17119
rect 24075 17085 24084 17119
rect 24032 17076 24084 17085
rect 24952 17076 25004 17128
rect 29644 17076 29696 17128
rect 33508 17076 33560 17128
rect 37280 17144 37332 17196
rect 38936 17144 38988 17196
rect 15292 17008 15344 17060
rect 17684 17008 17736 17060
rect 22560 17051 22612 17060
rect 22560 17017 22569 17051
rect 22569 17017 22603 17051
rect 22603 17017 22612 17051
rect 22560 17008 22612 17017
rect 16580 16940 16632 16992
rect 22192 16940 22244 16992
rect 27252 17008 27304 17060
rect 30196 17008 30248 17060
rect 35992 17051 36044 17060
rect 28172 16983 28224 16992
rect 28172 16949 28181 16983
rect 28181 16949 28215 16983
rect 28215 16949 28224 16983
rect 28172 16940 28224 16949
rect 34244 16983 34296 16992
rect 34244 16949 34253 16983
rect 34253 16949 34287 16983
rect 34287 16949 34296 16983
rect 34244 16940 34296 16949
rect 34888 16940 34940 16992
rect 35992 17017 36001 17051
rect 36001 17017 36035 17051
rect 36035 17017 36044 17051
rect 35992 17008 36044 17017
rect 36820 17051 36872 17060
rect 36820 17017 36829 17051
rect 36829 17017 36863 17051
rect 36863 17017 36872 17051
rect 36820 17008 36872 17017
rect 37832 17076 37884 17128
rect 38752 17119 38804 17128
rect 38752 17085 38761 17119
rect 38761 17085 38795 17119
rect 38795 17085 38804 17119
rect 38752 17076 38804 17085
rect 43996 17119 44048 17128
rect 43996 17085 44005 17119
rect 44005 17085 44039 17119
rect 44039 17085 44048 17119
rect 43996 17076 44048 17085
rect 44272 17119 44324 17128
rect 44272 17085 44281 17119
rect 44281 17085 44315 17119
rect 44315 17085 44324 17119
rect 44272 17076 44324 17085
rect 48872 17076 48924 17128
rect 50804 17076 50856 17128
rect 46204 17008 46256 17060
rect 39212 16940 39264 16992
rect 48504 16983 48556 16992
rect 48504 16949 48513 16983
rect 48513 16949 48547 16983
rect 48547 16949 48556 16983
rect 48504 16940 48556 16949
rect 49976 16983 50028 16992
rect 49976 16949 49985 16983
rect 49985 16949 50019 16983
rect 50019 16949 50028 16983
rect 49976 16940 50028 16949
rect 21344 16838 21396 16890
rect 21408 16838 21460 16890
rect 21472 16838 21524 16890
rect 21536 16838 21588 16890
rect 41707 16838 41759 16890
rect 41771 16838 41823 16890
rect 41835 16838 41887 16890
rect 41899 16838 41951 16890
rect 13820 16668 13872 16720
rect 14280 16668 14332 16720
rect 15292 16711 15344 16720
rect 15292 16677 15301 16711
rect 15301 16677 15335 16711
rect 15335 16677 15344 16711
rect 15292 16668 15344 16677
rect 11704 16600 11756 16652
rect 12532 16600 12584 16652
rect 18144 16736 18196 16788
rect 23940 16736 23992 16788
rect 33508 16736 33560 16788
rect 36820 16736 36872 16788
rect 39212 16779 39264 16788
rect 17684 16668 17736 16720
rect 22560 16668 22612 16720
rect 16672 16643 16724 16652
rect 16672 16609 16681 16643
rect 16681 16609 16715 16643
rect 16715 16609 16724 16643
rect 16672 16600 16724 16609
rect 16948 16643 17000 16652
rect 16948 16609 16957 16643
rect 16957 16609 16991 16643
rect 16991 16609 17000 16643
rect 16948 16600 17000 16609
rect 20076 16600 20128 16652
rect 29644 16668 29696 16720
rect 30196 16711 30248 16720
rect 30196 16677 30205 16711
rect 30205 16677 30239 16711
rect 30239 16677 30248 16711
rect 30196 16668 30248 16677
rect 39212 16745 39221 16779
rect 39221 16745 39255 16779
rect 39255 16745 39264 16779
rect 39212 16736 39264 16745
rect 46940 16736 46992 16788
rect 50804 16779 50856 16788
rect 50804 16745 50813 16779
rect 50813 16745 50847 16779
rect 50847 16745 50856 16779
rect 50804 16736 50856 16745
rect 29276 16600 29328 16652
rect 31392 16600 31444 16652
rect 34796 16600 34848 16652
rect 35164 16643 35216 16652
rect 35164 16609 35173 16643
rect 35173 16609 35207 16643
rect 35207 16609 35216 16643
rect 35164 16600 35216 16609
rect 37832 16643 37884 16652
rect 37832 16609 37841 16643
rect 37841 16609 37875 16643
rect 37875 16609 37884 16643
rect 37832 16600 37884 16609
rect 39212 16600 39264 16652
rect 40500 16643 40552 16652
rect 40500 16609 40509 16643
rect 40509 16609 40543 16643
rect 40543 16609 40552 16643
rect 40500 16600 40552 16609
rect 42892 16600 42944 16652
rect 43996 16600 44048 16652
rect 45928 16600 45980 16652
rect 48044 16600 48096 16652
rect 55312 16643 55364 16652
rect 55312 16609 55321 16643
rect 55321 16609 55355 16643
rect 55355 16609 55364 16643
rect 55312 16600 55364 16609
rect 55588 16643 55640 16652
rect 55588 16609 55597 16643
rect 55597 16609 55631 16643
rect 55631 16609 55640 16643
rect 55588 16600 55640 16609
rect 16488 16532 16540 16584
rect 18420 16532 18472 16584
rect 22744 16575 22796 16584
rect 22744 16541 22753 16575
rect 22753 16541 22787 16575
rect 22787 16541 22796 16575
rect 22744 16532 22796 16541
rect 23020 16575 23072 16584
rect 23020 16541 23029 16575
rect 23029 16541 23063 16575
rect 23063 16541 23072 16575
rect 23020 16532 23072 16541
rect 27988 16575 28040 16584
rect 27988 16541 27997 16575
rect 27997 16541 28031 16575
rect 28031 16541 28040 16575
rect 27988 16532 28040 16541
rect 32864 16532 32916 16584
rect 35256 16532 35308 16584
rect 35532 16532 35584 16584
rect 43720 16532 43772 16584
rect 46112 16575 46164 16584
rect 46112 16541 46121 16575
rect 46121 16541 46155 16575
rect 46155 16541 46164 16575
rect 46112 16532 46164 16541
rect 49700 16575 49752 16584
rect 49700 16541 49709 16575
rect 49709 16541 49743 16575
rect 49743 16541 49752 16575
rect 49700 16532 49752 16541
rect 57060 16532 57112 16584
rect 58440 16532 58492 16584
rect 18236 16396 18288 16448
rect 22928 16396 22980 16448
rect 28724 16396 28776 16448
rect 40592 16439 40644 16448
rect 40592 16405 40601 16439
rect 40601 16405 40635 16439
rect 40635 16405 40644 16439
rect 40592 16396 40644 16405
rect 43076 16396 43128 16448
rect 11163 16294 11215 16346
rect 11227 16294 11279 16346
rect 11291 16294 11343 16346
rect 11355 16294 11407 16346
rect 31526 16294 31578 16346
rect 31590 16294 31642 16346
rect 31654 16294 31706 16346
rect 31718 16294 31770 16346
rect 51888 16294 51940 16346
rect 51952 16294 52004 16346
rect 52016 16294 52068 16346
rect 52080 16294 52132 16346
rect 13084 16235 13136 16244
rect 13084 16201 13093 16235
rect 13093 16201 13127 16235
rect 13127 16201 13136 16235
rect 13084 16192 13136 16201
rect 18604 16192 18656 16244
rect 23664 16192 23716 16244
rect 12164 15988 12216 16040
rect 16304 16124 16356 16176
rect 25872 16192 25924 16244
rect 31392 16192 31444 16244
rect 34888 16192 34940 16244
rect 37372 16192 37424 16244
rect 39212 16235 39264 16244
rect 39212 16201 39221 16235
rect 39221 16201 39255 16235
rect 39255 16201 39264 16235
rect 39212 16192 39264 16201
rect 44272 16192 44324 16244
rect 48964 16192 49016 16244
rect 27896 16124 27948 16176
rect 15476 16056 15528 16108
rect 12716 15988 12768 16040
rect 14372 16031 14424 16040
rect 14372 15997 14381 16031
rect 14381 15997 14415 16031
rect 14415 15997 14424 16031
rect 14372 15988 14424 15997
rect 15200 15988 15252 16040
rect 18236 16031 18288 16040
rect 18236 15997 18245 16031
rect 18245 15997 18279 16031
rect 18279 15997 18288 16031
rect 18236 15988 18288 15997
rect 18328 16031 18380 16040
rect 18328 15997 18337 16031
rect 18337 15997 18371 16031
rect 18371 15997 18380 16031
rect 20628 16031 20680 16040
rect 18328 15988 18380 15997
rect 20628 15997 20637 16031
rect 20637 15997 20671 16031
rect 20671 15997 20680 16031
rect 20628 15988 20680 15997
rect 22284 16031 22336 16040
rect 2780 15920 2832 15972
rect 12348 15920 12400 15972
rect 940 15852 992 15904
rect 10140 15852 10192 15904
rect 15292 15920 15344 15972
rect 16580 15920 16632 15972
rect 17224 15920 17276 15972
rect 19524 15920 19576 15972
rect 22284 15997 22293 16031
rect 22293 15997 22327 16031
rect 22327 15997 22336 16031
rect 22284 15988 22336 15997
rect 21180 15963 21232 15972
rect 21180 15929 21189 15963
rect 21189 15929 21223 15963
rect 21223 15929 21232 15963
rect 21180 15920 21232 15929
rect 22192 15963 22244 15972
rect 22192 15929 22201 15963
rect 22201 15929 22235 15963
rect 22235 15929 22244 15963
rect 22192 15920 22244 15929
rect 27988 16099 28040 16108
rect 27988 16065 27997 16099
rect 27997 16065 28031 16099
rect 28031 16065 28040 16099
rect 27988 16056 28040 16065
rect 35256 16056 35308 16108
rect 37832 16056 37884 16108
rect 22836 15988 22888 16040
rect 24032 15988 24084 16040
rect 24860 15920 24912 15972
rect 29276 16031 29328 16040
rect 29276 15997 29285 16031
rect 29285 15997 29319 16031
rect 29319 15997 29328 16031
rect 29276 15988 29328 15997
rect 29552 16031 29604 16040
rect 29552 15997 29561 16031
rect 29561 15997 29595 16031
rect 29595 15997 29604 16031
rect 29552 15988 29604 15997
rect 33876 15988 33928 16040
rect 34888 16031 34940 16040
rect 34888 15997 34897 16031
rect 34897 15997 34931 16031
rect 34931 15997 34940 16031
rect 34888 15988 34940 15997
rect 35532 15988 35584 16040
rect 36544 16031 36596 16040
rect 36544 15997 36553 16031
rect 36553 15997 36587 16031
rect 36587 15997 36596 16031
rect 36544 15988 36596 15997
rect 38384 15988 38436 16040
rect 38936 16031 38988 16040
rect 38936 15997 38945 16031
rect 38945 15997 38979 16031
rect 38979 15997 38988 16031
rect 38936 15988 38988 15997
rect 28172 15920 28224 15972
rect 35348 15920 35400 15972
rect 38200 15920 38252 15972
rect 42064 15988 42116 16040
rect 46664 16056 46716 16108
rect 62304 16056 62356 16108
rect 43076 16031 43128 16040
rect 43076 15997 43085 16031
rect 43085 15997 43119 16031
rect 43119 15997 43128 16031
rect 43076 15988 43128 15997
rect 44088 15988 44140 16040
rect 44548 16031 44600 16040
rect 44548 15997 44557 16031
rect 44557 15997 44591 16031
rect 44591 15997 44600 16031
rect 44548 15988 44600 15997
rect 44732 15988 44784 16040
rect 46204 15988 46256 16040
rect 46940 15988 46992 16040
rect 48044 16031 48096 16040
rect 48044 15997 48053 16031
rect 48053 15997 48087 16031
rect 48087 15997 48096 16031
rect 48044 15988 48096 15997
rect 48320 16031 48372 16040
rect 48320 15997 48329 16031
rect 48329 15997 48363 16031
rect 48363 15997 48372 16031
rect 48320 15988 48372 15997
rect 57060 15988 57112 16040
rect 43628 15920 43680 15972
rect 44456 15963 44508 15972
rect 44456 15929 44465 15963
rect 44465 15929 44499 15963
rect 44499 15929 44508 15963
rect 44456 15920 44508 15929
rect 55128 15920 55180 15972
rect 27068 15852 27120 15904
rect 45192 15852 45244 15904
rect 55864 15895 55916 15904
rect 55864 15861 55873 15895
rect 55873 15861 55907 15895
rect 55907 15861 55916 15895
rect 55864 15852 55916 15861
rect 21344 15750 21396 15802
rect 21408 15750 21460 15802
rect 21472 15750 21524 15802
rect 21536 15750 21588 15802
rect 41707 15750 41759 15802
rect 41771 15750 41823 15802
rect 41835 15750 41887 15802
rect 41899 15750 41951 15802
rect 12348 15648 12400 15700
rect 27068 15648 27120 15700
rect 33876 15648 33928 15700
rect 36084 15648 36136 15700
rect 38384 15648 38436 15700
rect 4712 15580 4764 15632
rect 5448 15444 5500 15496
rect 6000 15512 6052 15564
rect 8116 15580 8168 15632
rect 17960 15580 18012 15632
rect 22008 15580 22060 15632
rect 22284 15580 22336 15632
rect 24952 15623 25004 15632
rect 24952 15589 24961 15623
rect 24961 15589 24995 15623
rect 24995 15589 25004 15623
rect 24952 15580 25004 15589
rect 28724 15623 28776 15632
rect 28724 15589 28733 15623
rect 28733 15589 28767 15623
rect 28767 15589 28776 15623
rect 28724 15580 28776 15589
rect 29552 15580 29604 15632
rect 35992 15580 36044 15632
rect 40592 15580 40644 15632
rect 43628 15623 43680 15632
rect 43628 15589 43637 15623
rect 43637 15589 43671 15623
rect 43671 15589 43680 15623
rect 43628 15580 43680 15589
rect 45192 15623 45244 15632
rect 45192 15589 45201 15623
rect 45201 15589 45235 15623
rect 45235 15589 45244 15623
rect 45192 15580 45244 15589
rect 46112 15580 46164 15632
rect 48504 15648 48556 15700
rect 48320 15580 48372 15632
rect 49976 15648 50028 15700
rect 49700 15623 49752 15632
rect 49700 15589 49709 15623
rect 49709 15589 49743 15623
rect 49743 15589 49752 15623
rect 49700 15580 49752 15589
rect 8576 15512 8628 15564
rect 10416 15512 10468 15564
rect 12164 15555 12216 15564
rect 12164 15521 12173 15555
rect 12173 15521 12207 15555
rect 12207 15521 12216 15555
rect 12164 15512 12216 15521
rect 13820 15555 13872 15564
rect 10324 15444 10376 15496
rect 13820 15521 13829 15555
rect 13829 15521 13863 15555
rect 13863 15521 13872 15555
rect 13820 15512 13872 15521
rect 15476 15555 15528 15564
rect 15476 15521 15485 15555
rect 15485 15521 15519 15555
rect 15519 15521 15528 15555
rect 15476 15512 15528 15521
rect 16672 15512 16724 15564
rect 17224 15555 17276 15564
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 19708 15512 19760 15564
rect 22836 15555 22888 15564
rect 22836 15521 22845 15555
rect 22845 15521 22879 15555
rect 22879 15521 22888 15555
rect 22836 15512 22888 15521
rect 23112 15512 23164 15564
rect 22376 15444 22428 15496
rect 23296 15487 23348 15496
rect 23296 15453 23305 15487
rect 23305 15453 23339 15487
rect 23339 15453 23348 15487
rect 23296 15444 23348 15453
rect 24492 15555 24544 15564
rect 24492 15521 24501 15555
rect 24501 15521 24535 15555
rect 24535 15521 24544 15555
rect 27068 15555 27120 15564
rect 24492 15512 24544 15521
rect 27068 15521 27077 15555
rect 27077 15521 27111 15555
rect 27111 15521 27120 15555
rect 27068 15512 27120 15521
rect 27528 15512 27580 15564
rect 28632 15512 28684 15564
rect 28816 15555 28868 15564
rect 28816 15521 28825 15555
rect 28825 15521 28859 15555
rect 28859 15521 28868 15555
rect 28816 15512 28868 15521
rect 36176 15512 36228 15564
rect 37740 15512 37792 15564
rect 38384 15555 38436 15564
rect 38384 15521 38393 15555
rect 38393 15521 38427 15555
rect 38427 15521 38436 15555
rect 38384 15512 38436 15521
rect 39028 15512 39080 15564
rect 44180 15512 44232 15564
rect 45284 15555 45336 15564
rect 45284 15521 45293 15555
rect 45293 15521 45327 15555
rect 45327 15521 45336 15555
rect 45284 15512 45336 15521
rect 46940 15512 46992 15564
rect 49240 15555 49292 15564
rect 49240 15521 49249 15555
rect 49249 15521 49283 15555
rect 49283 15521 49292 15555
rect 49240 15512 49292 15521
rect 49608 15512 49660 15564
rect 51632 15580 51684 15632
rect 52644 15580 52696 15632
rect 25504 15444 25556 15496
rect 32864 15487 32916 15496
rect 32864 15453 32873 15487
rect 32873 15453 32907 15487
rect 32907 15453 32916 15487
rect 32864 15444 32916 15453
rect 33140 15487 33192 15496
rect 33140 15453 33149 15487
rect 33149 15453 33183 15487
rect 33183 15453 33192 15487
rect 33140 15444 33192 15453
rect 36084 15487 36136 15496
rect 36084 15453 36093 15487
rect 36093 15453 36127 15487
rect 36127 15453 36136 15487
rect 36084 15444 36136 15453
rect 51540 15487 51592 15496
rect 51540 15453 51549 15487
rect 51549 15453 51583 15487
rect 51583 15453 51592 15487
rect 51540 15444 51592 15453
rect 15292 15376 15344 15428
rect 23664 15376 23716 15428
rect 27252 15419 27304 15428
rect 27252 15385 27261 15419
rect 27261 15385 27295 15419
rect 27295 15385 27304 15419
rect 27252 15376 27304 15385
rect 27896 15376 27948 15428
rect 33876 15376 33928 15428
rect 42064 15376 42116 15428
rect 43536 15376 43588 15428
rect 53288 15512 53340 15564
rect 58716 15580 58768 15632
rect 60372 15580 60424 15632
rect 52920 15487 52972 15496
rect 52920 15453 52929 15487
rect 52929 15453 52963 15487
rect 52963 15453 52972 15487
rect 52920 15444 52972 15453
rect 54668 15376 54720 15428
rect 55128 15376 55180 15428
rect 5356 15308 5408 15360
rect 7012 15308 7064 15360
rect 11060 15351 11112 15360
rect 11060 15317 11069 15351
rect 11069 15317 11103 15351
rect 11103 15317 11112 15351
rect 11060 15308 11112 15317
rect 12532 15351 12584 15360
rect 12532 15317 12541 15351
rect 12541 15317 12575 15351
rect 12575 15317 12584 15351
rect 12532 15308 12584 15317
rect 19616 15351 19668 15360
rect 19616 15317 19625 15351
rect 19625 15317 19659 15351
rect 19659 15317 19668 15351
rect 19616 15308 19668 15317
rect 27528 15308 27580 15360
rect 31116 15351 31168 15360
rect 31116 15317 31125 15351
rect 31125 15317 31159 15351
rect 31159 15317 31168 15351
rect 31116 15308 31168 15317
rect 33048 15308 33100 15360
rect 36544 15351 36596 15360
rect 36544 15317 36553 15351
rect 36553 15317 36587 15351
rect 36587 15317 36596 15351
rect 36544 15308 36596 15317
rect 38752 15351 38804 15360
rect 38752 15317 38761 15351
rect 38761 15317 38795 15351
rect 38795 15317 38804 15351
rect 38752 15308 38804 15317
rect 43720 15308 43772 15360
rect 44088 15308 44140 15360
rect 53288 15308 53340 15360
rect 54576 15308 54628 15360
rect 55496 15308 55548 15360
rect 11163 15206 11215 15258
rect 11227 15206 11279 15258
rect 11291 15206 11343 15258
rect 11355 15206 11407 15258
rect 31526 15206 31578 15258
rect 31590 15206 31642 15258
rect 31654 15206 31706 15258
rect 31718 15206 31770 15258
rect 51888 15206 51940 15258
rect 51952 15206 52004 15258
rect 52016 15206 52068 15258
rect 52080 15206 52132 15258
rect 8576 15147 8628 15156
rect 8576 15113 8585 15147
rect 8585 15113 8619 15147
rect 8619 15113 8628 15147
rect 8576 15104 8628 15113
rect 16304 15147 16356 15156
rect 16304 15113 16313 15147
rect 16313 15113 16347 15147
rect 16347 15113 16356 15147
rect 16304 15104 16356 15113
rect 16948 15104 17000 15156
rect 23020 15104 23072 15156
rect 25504 15147 25556 15156
rect 25504 15113 25513 15147
rect 25513 15113 25547 15147
rect 25547 15113 25556 15147
rect 25504 15104 25556 15113
rect 27896 15104 27948 15156
rect 28632 15104 28684 15156
rect 33048 15104 33100 15156
rect 33140 15104 33192 15156
rect 35164 15104 35216 15156
rect 37372 15104 37424 15156
rect 43536 15147 43588 15156
rect 43536 15113 43545 15147
rect 43545 15113 43579 15147
rect 43579 15113 43588 15147
rect 43536 15104 43588 15113
rect 44456 15104 44508 15156
rect 49608 15104 49660 15156
rect 53288 15147 53340 15156
rect 53288 15113 53297 15147
rect 53297 15113 53331 15147
rect 53331 15113 53340 15147
rect 53288 15104 53340 15113
rect 55588 15104 55640 15156
rect 12440 15036 12492 15088
rect 5448 14900 5500 14952
rect 6644 14900 6696 14952
rect 7104 14900 7156 14952
rect 7564 14900 7616 14952
rect 11704 14900 11756 14952
rect 12716 14943 12768 14952
rect 12716 14909 12725 14943
rect 12725 14909 12759 14943
rect 12759 14909 12768 14943
rect 12716 14900 12768 14909
rect 10968 14875 11020 14884
rect 10968 14841 10977 14875
rect 10977 14841 11011 14875
rect 11011 14841 11020 14875
rect 10968 14832 11020 14841
rect 12532 14832 12584 14884
rect 5632 14807 5684 14816
rect 5632 14773 5641 14807
rect 5641 14773 5675 14807
rect 5675 14773 5684 14807
rect 5632 14764 5684 14773
rect 10416 14764 10468 14816
rect 16488 14943 16540 14952
rect 16488 14909 16497 14943
rect 16497 14909 16531 14943
rect 16531 14909 16540 14943
rect 16488 14900 16540 14909
rect 16580 14943 16632 14952
rect 16580 14909 16589 14943
rect 16589 14909 16623 14943
rect 16623 14909 16632 14943
rect 16580 14900 16632 14909
rect 18420 14900 18472 14952
rect 18788 14943 18840 14952
rect 18788 14909 18797 14943
rect 18797 14909 18831 14943
rect 18831 14909 18840 14943
rect 18788 14900 18840 14909
rect 21180 14900 21232 14952
rect 22376 14900 22428 14952
rect 22744 14968 22796 15020
rect 23664 15011 23716 15020
rect 23664 14977 23673 15011
rect 23673 14977 23707 15011
rect 23707 14977 23716 15011
rect 23664 14968 23716 14977
rect 28172 15036 28224 15088
rect 23020 14900 23072 14952
rect 23296 14900 23348 14952
rect 25412 14943 25464 14952
rect 25412 14909 25421 14943
rect 25421 14909 25455 14943
rect 25455 14909 25464 14943
rect 25412 14900 25464 14909
rect 25504 14900 25556 14952
rect 27896 14900 27948 14952
rect 30932 14943 30984 14952
rect 30932 14909 30941 14943
rect 30941 14909 30975 14943
rect 30975 14909 30984 14943
rect 30932 14900 30984 14909
rect 32864 14900 32916 14952
rect 33324 14943 33376 14952
rect 33324 14909 33333 14943
rect 33333 14909 33367 14943
rect 33367 14909 33376 14943
rect 33324 14900 33376 14909
rect 36176 15036 36228 15088
rect 19432 14764 19484 14816
rect 19800 14764 19852 14816
rect 22928 14764 22980 14816
rect 27252 14832 27304 14884
rect 30748 14875 30800 14884
rect 30748 14841 30757 14875
rect 30757 14841 30791 14875
rect 30791 14841 30800 14875
rect 30748 14832 30800 14841
rect 33416 14875 33468 14884
rect 33416 14841 33425 14875
rect 33425 14841 33459 14875
rect 33459 14841 33468 14875
rect 33416 14832 33468 14841
rect 36084 14968 36136 15020
rect 37372 15011 37424 15020
rect 37372 14977 37381 15011
rect 37381 14977 37415 15011
rect 37415 14977 37424 15011
rect 37372 14968 37424 14977
rect 35348 14943 35400 14952
rect 35348 14909 35357 14943
rect 35357 14909 35391 14943
rect 35391 14909 35400 14943
rect 35348 14900 35400 14909
rect 36176 14900 36228 14952
rect 36636 14900 36688 14952
rect 24032 14764 24084 14816
rect 28816 14764 28868 14816
rect 30656 14764 30708 14816
rect 34612 14764 34664 14816
rect 38660 14900 38712 14952
rect 47032 14968 47084 15020
rect 50252 14968 50304 15020
rect 55312 14968 55364 15020
rect 41604 14900 41656 14952
rect 44364 14900 44416 14952
rect 45008 14900 45060 14952
rect 46664 14900 46716 14952
rect 40960 14832 41012 14884
rect 44732 14832 44784 14884
rect 53472 14900 53524 14952
rect 55036 14943 55088 14952
rect 55036 14909 55045 14943
rect 55045 14909 55079 14943
rect 55079 14909 55088 14943
rect 55036 14900 55088 14909
rect 55220 14943 55272 14952
rect 55220 14909 55229 14943
rect 55229 14909 55263 14943
rect 55263 14909 55272 14943
rect 55220 14900 55272 14909
rect 39120 14764 39172 14816
rect 43536 14764 43588 14816
rect 55864 14832 55916 14884
rect 46296 14764 46348 14816
rect 21344 14662 21396 14714
rect 21408 14662 21460 14714
rect 21472 14662 21524 14714
rect 21536 14662 21588 14714
rect 41707 14662 41759 14714
rect 41771 14662 41823 14714
rect 41835 14662 41887 14714
rect 41899 14662 41951 14714
rect 6000 14603 6052 14612
rect 6000 14569 6009 14603
rect 6009 14569 6043 14603
rect 6043 14569 6052 14603
rect 6000 14560 6052 14569
rect 6644 14560 6696 14612
rect 8116 14492 8168 14544
rect 10968 14560 11020 14612
rect 17960 14492 18012 14544
rect 20720 14492 20772 14544
rect 24860 14560 24912 14612
rect 7104 14467 7156 14476
rect 7104 14433 7113 14467
rect 7113 14433 7147 14467
rect 7147 14433 7156 14467
rect 10508 14467 10560 14476
rect 7104 14424 7156 14433
rect 5540 14356 5592 14408
rect 7380 14399 7432 14408
rect 7380 14365 7389 14399
rect 7389 14365 7423 14399
rect 7423 14365 7432 14399
rect 7380 14356 7432 14365
rect 10508 14433 10517 14467
rect 10517 14433 10551 14467
rect 10551 14433 10560 14467
rect 10508 14424 10560 14433
rect 11704 14399 11756 14408
rect 11704 14365 11713 14399
rect 11713 14365 11747 14399
rect 11747 14365 11756 14399
rect 11704 14356 11756 14365
rect 12992 14356 13044 14408
rect 15476 14424 15528 14476
rect 16672 14467 16724 14476
rect 16672 14433 16681 14467
rect 16681 14433 16715 14467
rect 16715 14433 16724 14467
rect 16672 14424 16724 14433
rect 19432 14467 19484 14476
rect 19432 14433 19441 14467
rect 19441 14433 19475 14467
rect 19475 14433 19484 14467
rect 19432 14424 19484 14433
rect 19524 14467 19576 14476
rect 19524 14433 19533 14467
rect 19533 14433 19567 14467
rect 19567 14433 19576 14467
rect 19524 14424 19576 14433
rect 17132 14356 17184 14408
rect 22376 14399 22428 14408
rect 22376 14365 22385 14399
rect 22385 14365 22419 14399
rect 22419 14365 22428 14399
rect 24492 14492 24544 14544
rect 22376 14356 22428 14365
rect 20168 14288 20220 14340
rect 24308 14467 24360 14476
rect 24308 14433 24317 14467
rect 24317 14433 24351 14467
rect 24351 14433 24360 14467
rect 24308 14424 24360 14433
rect 28908 14492 28960 14544
rect 24676 14467 24728 14476
rect 24676 14433 24685 14467
rect 24685 14433 24719 14467
rect 24719 14433 24728 14467
rect 24676 14424 24728 14433
rect 26608 14424 26660 14476
rect 26792 14424 26844 14476
rect 27896 14424 27948 14476
rect 29460 14467 29512 14476
rect 29460 14433 29469 14467
rect 29469 14433 29503 14467
rect 29503 14433 29512 14467
rect 29460 14424 29512 14433
rect 31116 14492 31168 14544
rect 39120 14560 39172 14612
rect 33048 14492 33100 14544
rect 30840 14467 30892 14476
rect 23020 14288 23072 14340
rect 3516 14220 3568 14272
rect 7288 14220 7340 14272
rect 14188 14220 14240 14272
rect 22376 14220 22428 14272
rect 28908 14288 28960 14340
rect 30840 14433 30849 14467
rect 30849 14433 30883 14467
rect 30883 14433 30892 14467
rect 33416 14492 33468 14544
rect 34244 14492 34296 14544
rect 37188 14492 37240 14544
rect 39028 14535 39080 14544
rect 39028 14501 39037 14535
rect 39037 14501 39071 14535
rect 39071 14501 39080 14535
rect 39028 14492 39080 14501
rect 30840 14424 30892 14433
rect 34612 14467 34664 14476
rect 34612 14433 34621 14467
rect 34621 14433 34655 14467
rect 34655 14433 34664 14467
rect 34612 14424 34664 14433
rect 35716 14424 35768 14476
rect 38568 14424 38620 14476
rect 41604 14560 41656 14612
rect 42064 14560 42116 14612
rect 43720 14492 43772 14544
rect 47216 14560 47268 14612
rect 51632 14603 51684 14612
rect 51632 14569 51641 14603
rect 51641 14569 51675 14603
rect 51675 14569 51684 14603
rect 51632 14560 51684 14569
rect 46664 14492 46716 14544
rect 52920 14535 52972 14544
rect 52920 14501 52929 14535
rect 52929 14501 52963 14535
rect 52963 14501 52972 14535
rect 52920 14492 52972 14501
rect 53472 14535 53524 14544
rect 53472 14501 53481 14535
rect 53481 14501 53515 14535
rect 53515 14501 53524 14535
rect 53472 14492 53524 14501
rect 56508 14492 56560 14544
rect 58716 14535 58768 14544
rect 58716 14501 58725 14535
rect 58725 14501 58759 14535
rect 58759 14501 58768 14535
rect 58716 14492 58768 14501
rect 43628 14467 43680 14476
rect 37648 14356 37700 14408
rect 38476 14356 38528 14408
rect 36084 14288 36136 14340
rect 38660 14288 38712 14340
rect 39396 14288 39448 14340
rect 39856 14356 39908 14408
rect 43628 14433 43637 14467
rect 43637 14433 43671 14467
rect 43671 14433 43680 14467
rect 43628 14424 43680 14433
rect 45928 14424 45980 14476
rect 46112 14424 46164 14476
rect 48044 14424 48096 14476
rect 50252 14467 50304 14476
rect 50252 14433 50261 14467
rect 50261 14433 50295 14467
rect 50295 14433 50304 14467
rect 50252 14424 50304 14433
rect 53012 14467 53064 14476
rect 53012 14433 53021 14467
rect 53021 14433 53055 14467
rect 53055 14433 53064 14467
rect 53012 14424 53064 14433
rect 55312 14424 55364 14476
rect 44456 14356 44508 14408
rect 46572 14356 46624 14408
rect 52184 14356 52236 14408
rect 54852 14399 54904 14408
rect 54852 14365 54861 14399
rect 54861 14365 54895 14399
rect 54895 14365 54904 14399
rect 54852 14356 54904 14365
rect 56416 14356 56468 14408
rect 57336 14399 57388 14408
rect 57336 14365 57345 14399
rect 57345 14365 57379 14399
rect 57379 14365 57388 14399
rect 57336 14356 57388 14365
rect 40776 14288 40828 14340
rect 30932 14220 30984 14272
rect 32496 14220 32548 14272
rect 34796 14263 34848 14272
rect 34796 14229 34805 14263
rect 34805 14229 34839 14263
rect 34839 14229 34848 14263
rect 34796 14220 34848 14229
rect 34888 14220 34940 14272
rect 39120 14220 39172 14272
rect 45468 14220 45520 14272
rect 52736 14263 52788 14272
rect 52736 14229 52745 14263
rect 52745 14229 52779 14263
rect 52779 14229 52788 14263
rect 52736 14220 52788 14229
rect 11163 14118 11215 14170
rect 11227 14118 11279 14170
rect 11291 14118 11343 14170
rect 11355 14118 11407 14170
rect 31526 14118 31578 14170
rect 31590 14118 31642 14170
rect 31654 14118 31706 14170
rect 31718 14118 31770 14170
rect 51888 14118 51940 14170
rect 51952 14118 52004 14170
rect 52016 14118 52068 14170
rect 52080 14118 52132 14170
rect 5264 14016 5316 14068
rect 11060 14016 11112 14068
rect 12348 14016 12400 14068
rect 12716 14016 12768 14068
rect 12992 14016 13044 14068
rect 22468 14059 22520 14068
rect 5264 13855 5316 13864
rect 5264 13821 5273 13855
rect 5273 13821 5307 13855
rect 5307 13821 5316 13855
rect 5264 13812 5316 13821
rect 5632 13880 5684 13932
rect 7196 13948 7248 14000
rect 7288 13948 7340 14000
rect 22468 14025 22477 14059
rect 22477 14025 22511 14059
rect 22511 14025 22520 14059
rect 22468 14016 22520 14025
rect 24308 14016 24360 14068
rect 24124 13948 24176 14000
rect 29276 14016 29328 14068
rect 29460 14016 29512 14068
rect 33324 14016 33376 14068
rect 38568 14016 38620 14068
rect 44180 14016 44232 14068
rect 44364 14016 44416 14068
rect 46112 14059 46164 14068
rect 46112 14025 46121 14059
rect 46121 14025 46155 14059
rect 46155 14025 46164 14059
rect 46112 14016 46164 14025
rect 46572 14059 46624 14068
rect 46572 14025 46581 14059
rect 46581 14025 46615 14059
rect 46615 14025 46624 14059
rect 46572 14016 46624 14025
rect 52184 14059 52236 14068
rect 52184 14025 52193 14059
rect 52193 14025 52227 14059
rect 52227 14025 52236 14059
rect 52184 14016 52236 14025
rect 52736 14016 52788 14068
rect 55036 14016 55088 14068
rect 7380 13880 7432 13932
rect 7564 13923 7616 13932
rect 7564 13889 7573 13923
rect 7573 13889 7607 13923
rect 7607 13889 7616 13923
rect 7564 13880 7616 13889
rect 12348 13880 12400 13932
rect 18144 13923 18196 13932
rect 18144 13889 18153 13923
rect 18153 13889 18187 13923
rect 18187 13889 18196 13923
rect 18144 13880 18196 13889
rect 18420 13880 18472 13932
rect 23020 13880 23072 13932
rect 25872 13923 25924 13932
rect 5816 13812 5868 13864
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 8300 13812 8352 13864
rect 11060 13855 11112 13864
rect 11060 13821 11069 13855
rect 11069 13821 11103 13855
rect 11103 13821 11112 13855
rect 11060 13812 11112 13821
rect 11520 13855 11572 13864
rect 10324 13787 10376 13796
rect 10324 13753 10333 13787
rect 10333 13753 10367 13787
rect 10367 13753 10376 13787
rect 10324 13744 10376 13753
rect 11520 13821 11529 13855
rect 11529 13821 11563 13855
rect 11563 13821 11572 13855
rect 11520 13812 11572 13821
rect 12716 13855 12768 13864
rect 12716 13821 12725 13855
rect 12725 13821 12759 13855
rect 12759 13821 12768 13855
rect 12716 13812 12768 13821
rect 13728 13812 13780 13864
rect 18236 13855 18288 13864
rect 18236 13821 18245 13855
rect 18245 13821 18279 13855
rect 18279 13821 18288 13855
rect 18236 13812 18288 13821
rect 20904 13812 20956 13864
rect 22100 13855 22152 13864
rect 22100 13821 22109 13855
rect 22109 13821 22143 13855
rect 22143 13821 22152 13855
rect 22284 13855 22336 13864
rect 22100 13812 22152 13821
rect 22284 13821 22293 13855
rect 22293 13821 22327 13855
rect 22327 13821 22336 13855
rect 22284 13812 22336 13821
rect 22376 13812 22428 13864
rect 25872 13889 25881 13923
rect 25881 13889 25915 13923
rect 25915 13889 25924 13923
rect 25872 13880 25924 13889
rect 11704 13744 11756 13796
rect 12532 13744 12584 13796
rect 14188 13787 14240 13796
rect 14188 13753 14197 13787
rect 14197 13753 14231 13787
rect 14231 13753 14240 13787
rect 14188 13744 14240 13753
rect 15384 13744 15436 13796
rect 18328 13744 18380 13796
rect 3332 13676 3384 13728
rect 21732 13676 21784 13728
rect 26608 13880 26660 13932
rect 29276 13880 29328 13932
rect 37372 13948 37424 14000
rect 37648 13948 37700 14000
rect 43720 13948 43772 14000
rect 26148 13855 26200 13864
rect 26148 13821 26157 13855
rect 26157 13821 26191 13855
rect 26191 13821 26200 13855
rect 26148 13812 26200 13821
rect 30472 13855 30524 13864
rect 30472 13821 30481 13855
rect 30481 13821 30515 13855
rect 30515 13821 30524 13855
rect 30472 13812 30524 13821
rect 30748 13812 30800 13864
rect 27068 13744 27120 13796
rect 30288 13744 30340 13796
rect 32864 13812 32916 13864
rect 36820 13855 36872 13864
rect 36820 13821 36829 13855
rect 36829 13821 36863 13855
rect 36863 13821 36872 13855
rect 36820 13812 36872 13821
rect 39120 13880 39172 13932
rect 47400 13880 47452 13932
rect 48228 13880 48280 13932
rect 38660 13812 38712 13864
rect 38844 13855 38896 13864
rect 38844 13821 38853 13855
rect 38853 13821 38887 13855
rect 38887 13821 38896 13855
rect 38844 13812 38896 13821
rect 39396 13855 39448 13864
rect 35164 13744 35216 13796
rect 36176 13787 36228 13796
rect 36176 13753 36185 13787
rect 36185 13753 36219 13787
rect 36219 13753 36228 13787
rect 36176 13744 36228 13753
rect 38200 13787 38252 13796
rect 38200 13753 38209 13787
rect 38209 13753 38243 13787
rect 38243 13753 38252 13787
rect 38200 13744 38252 13753
rect 31116 13676 31168 13728
rect 37372 13676 37424 13728
rect 38476 13676 38528 13728
rect 39396 13821 39405 13855
rect 39405 13821 39439 13855
rect 39439 13821 39448 13855
rect 39396 13812 39448 13821
rect 39856 13812 39908 13864
rect 44088 13812 44140 13864
rect 44732 13855 44784 13864
rect 44732 13821 44741 13855
rect 44741 13821 44775 13855
rect 44775 13821 44784 13855
rect 44732 13812 44784 13821
rect 44916 13812 44968 13864
rect 45652 13812 45704 13864
rect 46388 13855 46440 13864
rect 46388 13821 46397 13855
rect 46397 13821 46431 13855
rect 46431 13821 46440 13855
rect 46388 13812 46440 13821
rect 47032 13812 47084 13864
rect 46296 13787 46348 13796
rect 46296 13753 46305 13787
rect 46305 13753 46339 13787
rect 46339 13753 46348 13787
rect 46296 13744 46348 13753
rect 47216 13744 47268 13796
rect 51540 13880 51592 13932
rect 54852 13880 54904 13932
rect 52552 13812 52604 13864
rect 54024 13855 54076 13864
rect 54024 13821 54033 13855
rect 54033 13821 54067 13855
rect 54067 13821 54076 13855
rect 54024 13812 54076 13821
rect 54576 13812 54628 13864
rect 55496 13855 55548 13864
rect 55496 13821 55505 13855
rect 55505 13821 55539 13855
rect 55539 13821 55548 13855
rect 55496 13812 55548 13821
rect 57336 13880 57388 13932
rect 53564 13744 53616 13796
rect 53932 13787 53984 13796
rect 53932 13753 53941 13787
rect 53941 13753 53975 13787
rect 53975 13753 53984 13787
rect 53932 13744 53984 13753
rect 46204 13676 46256 13728
rect 48136 13676 48188 13728
rect 50068 13676 50120 13728
rect 21344 13574 21396 13626
rect 21408 13574 21460 13626
rect 21472 13574 21524 13626
rect 21536 13574 21588 13626
rect 41707 13574 41759 13626
rect 41771 13574 41823 13626
rect 41835 13574 41887 13626
rect 41899 13574 41951 13626
rect 4068 13472 4120 13524
rect 18880 13472 18932 13524
rect 19064 13472 19116 13524
rect 22652 13472 22704 13524
rect 5356 13447 5408 13456
rect 5356 13413 5365 13447
rect 5365 13413 5399 13447
rect 5399 13413 5408 13447
rect 5356 13404 5408 13413
rect 10416 13447 10468 13456
rect 10416 13413 10425 13447
rect 10425 13413 10459 13447
rect 10459 13413 10468 13447
rect 10416 13404 10468 13413
rect 15384 13404 15436 13456
rect 17132 13447 17184 13456
rect 17132 13413 17141 13447
rect 17141 13413 17175 13447
rect 17175 13413 17184 13447
rect 17132 13404 17184 13413
rect 18788 13404 18840 13456
rect 20904 13447 20956 13456
rect 20904 13413 20913 13447
rect 20913 13413 20947 13447
rect 20947 13413 20956 13447
rect 20904 13404 20956 13413
rect 24400 13472 24452 13524
rect 26792 13472 26844 13524
rect 26884 13472 26936 13524
rect 42892 13515 42944 13524
rect 5264 13379 5316 13388
rect 5264 13345 5273 13379
rect 5273 13345 5307 13379
rect 5307 13345 5316 13379
rect 5264 13336 5316 13345
rect 5448 13379 5500 13388
rect 5448 13345 5457 13379
rect 5457 13345 5491 13379
rect 5491 13345 5500 13379
rect 9772 13379 9824 13388
rect 5448 13336 5500 13345
rect 9772 13345 9781 13379
rect 9781 13345 9815 13379
rect 9815 13345 9824 13379
rect 9772 13336 9824 13345
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 11060 13268 11112 13320
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 12256 13336 12308 13388
rect 14648 13336 14700 13388
rect 15292 13379 15344 13388
rect 15292 13345 15301 13379
rect 15301 13345 15335 13379
rect 15335 13345 15344 13379
rect 15292 13336 15344 13345
rect 17040 13336 17092 13388
rect 17960 13379 18012 13388
rect 17960 13345 17969 13379
rect 17969 13345 18003 13379
rect 18003 13345 18012 13379
rect 17960 13336 18012 13345
rect 19524 13336 19576 13388
rect 19800 13379 19852 13388
rect 19800 13345 19809 13379
rect 19809 13345 19843 13379
rect 19843 13345 19852 13379
rect 19800 13336 19852 13345
rect 21180 13336 21232 13388
rect 21732 13379 21784 13388
rect 12348 13268 12400 13320
rect 13268 13268 13320 13320
rect 13452 13311 13504 13320
rect 13452 13277 13461 13311
rect 13461 13277 13495 13311
rect 13495 13277 13504 13311
rect 13452 13268 13504 13277
rect 12900 13200 12952 13252
rect 5540 13132 5592 13184
rect 10140 13132 10192 13184
rect 13636 13200 13688 13252
rect 13084 13132 13136 13184
rect 21732 13345 21741 13379
rect 21741 13345 21775 13379
rect 21775 13345 21784 13379
rect 21732 13336 21784 13345
rect 23020 13336 23072 13388
rect 24216 13336 24268 13388
rect 25228 13336 25280 13388
rect 27068 13379 27120 13388
rect 27068 13345 27077 13379
rect 27077 13345 27111 13379
rect 27111 13345 27120 13379
rect 27068 13336 27120 13345
rect 27344 13379 27396 13388
rect 27344 13345 27353 13379
rect 27353 13345 27387 13379
rect 27387 13345 27396 13379
rect 27344 13336 27396 13345
rect 27988 13336 28040 13388
rect 30380 13379 30432 13388
rect 30380 13345 30389 13379
rect 30389 13345 30423 13379
rect 30423 13345 30432 13379
rect 30380 13336 30432 13345
rect 30748 13379 30800 13388
rect 17224 13200 17276 13252
rect 28264 13268 28316 13320
rect 28448 13268 28500 13320
rect 30748 13345 30757 13379
rect 30757 13345 30791 13379
rect 30791 13345 30800 13379
rect 30748 13336 30800 13345
rect 32036 13404 32088 13456
rect 34888 13404 34940 13456
rect 36820 13404 36872 13456
rect 37740 13447 37792 13456
rect 37740 13413 37749 13447
rect 37749 13413 37783 13447
rect 37783 13413 37792 13447
rect 37740 13404 37792 13413
rect 42892 13481 42901 13515
rect 42901 13481 42935 13515
rect 42935 13481 42944 13515
rect 42892 13472 42944 13481
rect 53932 13472 53984 13524
rect 41328 13404 41380 13456
rect 42064 13404 42116 13456
rect 45284 13404 45336 13456
rect 49240 13404 49292 13456
rect 53012 13404 53064 13456
rect 54668 13447 54720 13456
rect 54668 13413 54677 13447
rect 54677 13413 54711 13447
rect 54711 13413 54720 13447
rect 54668 13404 54720 13413
rect 32404 13379 32456 13388
rect 32404 13345 32413 13379
rect 32413 13345 32447 13379
rect 32447 13345 32456 13379
rect 32404 13336 32456 13345
rect 33876 13268 33928 13320
rect 26240 13200 26292 13252
rect 22836 13132 22888 13184
rect 24308 13175 24360 13184
rect 24308 13141 24317 13175
rect 24317 13141 24351 13175
rect 24351 13141 24360 13175
rect 24308 13132 24360 13141
rect 25780 13132 25832 13184
rect 30104 13200 30156 13252
rect 30472 13200 30524 13252
rect 31116 13200 31168 13252
rect 35164 13336 35216 13388
rect 36176 13379 36228 13388
rect 36176 13345 36185 13379
rect 36185 13345 36219 13379
rect 36219 13345 36228 13379
rect 36176 13336 36228 13345
rect 38384 13379 38436 13388
rect 38384 13345 38393 13379
rect 38393 13345 38427 13379
rect 38427 13345 38436 13379
rect 38384 13336 38436 13345
rect 38476 13379 38528 13388
rect 38476 13345 38485 13379
rect 38485 13345 38519 13379
rect 38519 13345 38528 13379
rect 38476 13336 38528 13345
rect 35072 13268 35124 13320
rect 28724 13132 28776 13184
rect 30288 13132 30340 13184
rect 30932 13132 30984 13184
rect 36360 13200 36412 13252
rect 39396 13336 39448 13388
rect 41604 13336 41656 13388
rect 43076 13379 43128 13388
rect 43076 13345 43085 13379
rect 43085 13345 43119 13379
rect 43119 13345 43128 13379
rect 43076 13336 43128 13345
rect 43168 13336 43220 13388
rect 45744 13336 45796 13388
rect 46112 13336 46164 13388
rect 47124 13336 47176 13388
rect 47584 13336 47636 13388
rect 44364 13268 44416 13320
rect 44732 13268 44784 13320
rect 45652 13311 45704 13320
rect 45652 13277 45661 13311
rect 45661 13277 45695 13311
rect 45695 13277 45704 13311
rect 45652 13268 45704 13277
rect 45836 13268 45888 13320
rect 46480 13200 46532 13252
rect 46940 13243 46992 13252
rect 46940 13209 46949 13243
rect 46949 13209 46983 13243
rect 46983 13209 46992 13243
rect 46940 13200 46992 13209
rect 47400 13311 47452 13320
rect 47400 13277 47409 13311
rect 47409 13277 47443 13311
rect 47443 13277 47452 13311
rect 47400 13268 47452 13277
rect 48136 13336 48188 13388
rect 49608 13379 49660 13388
rect 49608 13345 49617 13379
rect 49617 13345 49651 13379
rect 49651 13345 49660 13379
rect 49608 13336 49660 13345
rect 49976 13379 50028 13388
rect 49976 13345 49985 13379
rect 49985 13345 50019 13379
rect 50019 13345 50028 13379
rect 49976 13336 50028 13345
rect 51172 13379 51224 13388
rect 51172 13345 51181 13379
rect 51181 13345 51215 13379
rect 51215 13345 51224 13379
rect 51172 13336 51224 13345
rect 53104 13379 53156 13388
rect 53104 13345 53113 13379
rect 53113 13345 53147 13379
rect 53147 13345 53156 13379
rect 53104 13336 53156 13345
rect 53380 13336 53432 13388
rect 56508 13336 56560 13388
rect 48228 13268 48280 13320
rect 50068 13311 50120 13320
rect 50068 13277 50077 13311
rect 50077 13277 50111 13311
rect 50111 13277 50120 13311
rect 50068 13268 50120 13277
rect 50620 13268 50672 13320
rect 51632 13311 51684 13320
rect 51632 13277 51641 13311
rect 51641 13277 51675 13311
rect 51675 13277 51684 13311
rect 51632 13268 51684 13277
rect 53196 13311 53248 13320
rect 53196 13277 53205 13311
rect 53205 13277 53239 13311
rect 53239 13277 53248 13311
rect 53196 13268 53248 13277
rect 53564 13311 53616 13320
rect 53564 13277 53573 13311
rect 53573 13277 53607 13311
rect 53607 13277 53616 13311
rect 53564 13268 53616 13277
rect 33692 13175 33744 13184
rect 33692 13141 33701 13175
rect 33701 13141 33735 13175
rect 33735 13141 33744 13175
rect 33692 13132 33744 13141
rect 33784 13132 33836 13184
rect 34244 13132 34296 13184
rect 40500 13132 40552 13184
rect 41420 13132 41472 13184
rect 45928 13132 45980 13184
rect 46664 13132 46716 13184
rect 11163 13030 11215 13082
rect 11227 13030 11279 13082
rect 11291 13030 11343 13082
rect 11355 13030 11407 13082
rect 31526 13030 31578 13082
rect 31590 13030 31642 13082
rect 31654 13030 31706 13082
rect 31718 13030 31770 13082
rect 51888 13030 51940 13082
rect 51952 13030 52004 13082
rect 52016 13030 52068 13082
rect 52080 13030 52132 13082
rect 5448 12928 5500 12980
rect 3056 12860 3108 12912
rect 5632 12724 5684 12776
rect 8944 12860 8996 12912
rect 12624 12928 12676 12980
rect 17224 12928 17276 12980
rect 18144 12928 18196 12980
rect 20352 12928 20404 12980
rect 7288 12792 7340 12844
rect 8300 12792 8352 12844
rect 6460 12724 6512 12776
rect 7472 12724 7524 12776
rect 7012 12656 7064 12708
rect 6552 12588 6604 12640
rect 9220 12767 9272 12776
rect 9220 12733 9229 12767
rect 9229 12733 9263 12767
rect 9263 12733 9272 12767
rect 9220 12724 9272 12733
rect 9312 12724 9364 12776
rect 11060 12767 11112 12776
rect 11060 12733 11069 12767
rect 11069 12733 11103 12767
rect 11103 12733 11112 12767
rect 11060 12724 11112 12733
rect 11520 12767 11572 12776
rect 11244 12656 11296 12708
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 11980 12724 12032 12776
rect 13268 12792 13320 12844
rect 13084 12767 13136 12776
rect 13084 12733 13093 12767
rect 13093 12733 13127 12767
rect 13127 12733 13136 12767
rect 13084 12724 13136 12733
rect 13360 12724 13412 12776
rect 14004 12724 14056 12776
rect 15752 12767 15804 12776
rect 15752 12733 15761 12767
rect 15761 12733 15795 12767
rect 15795 12733 15804 12767
rect 15752 12724 15804 12733
rect 17592 12860 17644 12912
rect 19616 12860 19668 12912
rect 20444 12860 20496 12912
rect 24308 12928 24360 12980
rect 30840 12928 30892 12980
rect 32036 12971 32088 12980
rect 16672 12724 16724 12776
rect 17592 12724 17644 12776
rect 20628 12792 20680 12844
rect 25780 12860 25832 12912
rect 26148 12860 26200 12912
rect 26240 12860 26292 12912
rect 32036 12937 32045 12971
rect 32045 12937 32079 12971
rect 32079 12937 32088 12971
rect 32036 12928 32088 12937
rect 40592 12928 40644 12980
rect 40776 12971 40828 12980
rect 40776 12937 40785 12971
rect 40785 12937 40819 12971
rect 40819 12937 40828 12971
rect 40776 12928 40828 12937
rect 43076 12928 43128 12980
rect 46112 12928 46164 12980
rect 46388 12928 46440 12980
rect 49608 12928 49660 12980
rect 54024 12928 54076 12980
rect 55220 12928 55272 12980
rect 20076 12724 20128 12776
rect 20260 12724 20312 12776
rect 20812 12767 20864 12776
rect 20812 12733 20821 12767
rect 20821 12733 20855 12767
rect 20855 12733 20864 12767
rect 20812 12724 20864 12733
rect 15200 12656 15252 12708
rect 12532 12588 12584 12640
rect 14648 12631 14700 12640
rect 14648 12597 14657 12631
rect 14657 12597 14691 12631
rect 14691 12597 14700 12631
rect 14648 12588 14700 12597
rect 16580 12588 16632 12640
rect 18788 12656 18840 12708
rect 18880 12656 18932 12708
rect 19432 12656 19484 12708
rect 19340 12588 19392 12640
rect 22100 12767 22152 12776
rect 22100 12733 22109 12767
rect 22109 12733 22143 12767
rect 22143 12733 22152 12767
rect 23664 12767 23716 12776
rect 22100 12724 22152 12733
rect 23664 12733 23673 12767
rect 23673 12733 23707 12767
rect 23707 12733 23716 12767
rect 23664 12724 23716 12733
rect 23940 12724 23992 12776
rect 26608 12792 26660 12844
rect 28448 12792 28500 12844
rect 26332 12656 26384 12708
rect 24400 12588 24452 12640
rect 26792 12724 26844 12776
rect 27712 12724 27764 12776
rect 28540 12724 28592 12776
rect 29368 12656 29420 12708
rect 27620 12588 27672 12640
rect 27896 12588 27948 12640
rect 30656 12724 30708 12776
rect 34428 12792 34480 12844
rect 32588 12767 32640 12776
rect 32588 12733 32597 12767
rect 32597 12733 32631 12767
rect 32631 12733 32640 12767
rect 32588 12724 32640 12733
rect 32956 12767 33008 12776
rect 32956 12733 32965 12767
rect 32965 12733 32999 12767
rect 32999 12733 33008 12767
rect 32956 12724 33008 12733
rect 38384 12792 38436 12844
rect 40500 12835 40552 12844
rect 40500 12801 40509 12835
rect 40509 12801 40543 12835
rect 40543 12801 40552 12835
rect 40500 12792 40552 12801
rect 43168 12792 43220 12844
rect 45100 12792 45152 12844
rect 47032 12860 47084 12912
rect 48228 12860 48280 12912
rect 47216 12835 47268 12844
rect 47216 12801 47225 12835
rect 47225 12801 47259 12835
rect 47259 12801 47268 12835
rect 47216 12792 47268 12801
rect 53196 12835 53248 12844
rect 53196 12801 53205 12835
rect 53205 12801 53239 12835
rect 53239 12801 53248 12835
rect 53196 12792 53248 12801
rect 53564 12792 53616 12844
rect 55036 12792 55088 12844
rect 56416 12792 56468 12844
rect 35900 12724 35952 12776
rect 36084 12767 36136 12776
rect 36084 12733 36093 12767
rect 36093 12733 36127 12767
rect 36127 12733 36136 12767
rect 36084 12724 36136 12733
rect 36176 12767 36228 12776
rect 36176 12733 36205 12767
rect 36205 12733 36228 12767
rect 36176 12724 36228 12733
rect 29644 12588 29696 12640
rect 33508 12656 33560 12708
rect 36544 12724 36596 12776
rect 37464 12767 37516 12776
rect 37464 12733 37473 12767
rect 37473 12733 37507 12767
rect 37507 12733 37516 12767
rect 37464 12724 37516 12733
rect 35164 12631 35216 12640
rect 35164 12597 35173 12631
rect 35173 12597 35207 12631
rect 35207 12597 35216 12631
rect 35164 12588 35216 12597
rect 36176 12588 36228 12640
rect 38844 12724 38896 12776
rect 40684 12724 40736 12776
rect 44364 12767 44416 12776
rect 43444 12656 43496 12708
rect 44364 12733 44373 12767
rect 44373 12733 44407 12767
rect 44407 12733 44416 12767
rect 44364 12724 44416 12733
rect 45376 12767 45428 12776
rect 45376 12733 45385 12767
rect 45385 12733 45419 12767
rect 45419 12733 45428 12767
rect 45376 12724 45428 12733
rect 47032 12724 47084 12776
rect 48136 12767 48188 12776
rect 48136 12733 48145 12767
rect 48145 12733 48179 12767
rect 48179 12733 48188 12767
rect 48136 12724 48188 12733
rect 50252 12767 50304 12776
rect 50252 12733 50261 12767
rect 50261 12733 50295 12767
rect 50295 12733 50304 12767
rect 50252 12724 50304 12733
rect 51080 12724 51132 12776
rect 51632 12724 51684 12776
rect 55312 12767 55364 12776
rect 48044 12656 48096 12708
rect 50068 12656 50120 12708
rect 50896 12656 50948 12708
rect 52736 12656 52788 12708
rect 55312 12733 55321 12767
rect 55321 12733 55355 12767
rect 55355 12733 55364 12767
rect 55312 12724 55364 12733
rect 55772 12767 55824 12776
rect 55772 12733 55781 12767
rect 55781 12733 55815 12767
rect 55815 12733 55824 12767
rect 55772 12724 55824 12733
rect 58440 12724 58492 12776
rect 56140 12656 56192 12708
rect 59728 12631 59780 12640
rect 59728 12597 59737 12631
rect 59737 12597 59771 12631
rect 59771 12597 59780 12631
rect 59728 12588 59780 12597
rect 21344 12486 21396 12538
rect 21408 12486 21460 12538
rect 21472 12486 21524 12538
rect 21536 12486 21588 12538
rect 41707 12486 41759 12538
rect 41771 12486 41823 12538
rect 41835 12486 41887 12538
rect 41899 12486 41951 12538
rect 2780 12384 2832 12436
rect 9864 12384 9916 12436
rect 5816 12316 5868 12368
rect 6460 12316 6512 12368
rect 6368 12291 6420 12300
rect 5632 12180 5684 12232
rect 6368 12257 6377 12291
rect 6377 12257 6411 12291
rect 6411 12257 6420 12291
rect 6368 12248 6420 12257
rect 7472 12291 7524 12300
rect 7472 12257 7481 12291
rect 7481 12257 7515 12291
rect 7515 12257 7524 12291
rect 7472 12248 7524 12257
rect 6828 12180 6880 12232
rect 9312 12316 9364 12368
rect 11152 12384 11204 12436
rect 11428 12316 11480 12368
rect 10784 12248 10836 12300
rect 11520 12291 11572 12300
rect 11520 12257 11529 12291
rect 11529 12257 11563 12291
rect 11563 12257 11572 12291
rect 11520 12248 11572 12257
rect 11888 12291 11940 12300
rect 11888 12257 11897 12291
rect 11897 12257 11931 12291
rect 11931 12257 11940 12291
rect 11888 12248 11940 12257
rect 12348 12316 12400 12368
rect 18880 12384 18932 12436
rect 16120 12316 16172 12368
rect 19340 12316 19392 12368
rect 15016 12248 15068 12300
rect 16672 12248 16724 12300
rect 17592 12291 17644 12300
rect 17592 12257 17601 12291
rect 17601 12257 17635 12291
rect 17635 12257 17644 12291
rect 17592 12248 17644 12257
rect 17776 12248 17828 12300
rect 19708 12316 19760 12368
rect 21640 12316 21692 12368
rect 19800 12291 19852 12300
rect 19800 12257 19809 12291
rect 19809 12257 19843 12291
rect 19843 12257 19852 12291
rect 19800 12248 19852 12257
rect 21732 12291 21784 12300
rect 7932 12180 7984 12232
rect 10968 12180 11020 12232
rect 11428 12223 11480 12232
rect 11428 12189 11437 12223
rect 11437 12189 11471 12223
rect 11471 12189 11480 12223
rect 11428 12180 11480 12189
rect 12900 12223 12952 12232
rect 12900 12189 12909 12223
rect 12909 12189 12943 12223
rect 12943 12189 12952 12223
rect 12900 12180 12952 12189
rect 7104 12112 7156 12164
rect 7564 12112 7616 12164
rect 13084 12112 13136 12164
rect 16396 12112 16448 12164
rect 21088 12180 21140 12232
rect 21732 12257 21741 12291
rect 21741 12257 21775 12291
rect 21775 12257 21784 12291
rect 21732 12248 21784 12257
rect 22284 12384 22336 12436
rect 23848 12384 23900 12436
rect 24400 12384 24452 12436
rect 30012 12384 30064 12436
rect 41420 12384 41472 12436
rect 23572 12248 23624 12300
rect 24124 12291 24176 12300
rect 24124 12257 24133 12291
rect 24133 12257 24167 12291
rect 24167 12257 24176 12291
rect 24124 12248 24176 12257
rect 25228 12248 25280 12300
rect 25412 12248 25464 12300
rect 28724 12291 28776 12300
rect 23480 12180 23532 12232
rect 24308 12180 24360 12232
rect 28724 12257 28733 12291
rect 28733 12257 28767 12291
rect 28767 12257 28776 12291
rect 28724 12248 28776 12257
rect 28816 12248 28868 12300
rect 29644 12316 29696 12368
rect 30104 12316 30156 12368
rect 30196 12248 30248 12300
rect 30748 12359 30800 12368
rect 30748 12325 30757 12359
rect 30757 12325 30791 12359
rect 30791 12325 30800 12359
rect 30748 12316 30800 12325
rect 31024 12316 31076 12368
rect 32404 12316 32456 12368
rect 28080 12223 28132 12232
rect 28080 12189 28089 12223
rect 28089 12189 28123 12223
rect 28123 12189 28132 12223
rect 28080 12180 28132 12189
rect 21548 12112 21600 12164
rect 22008 12112 22060 12164
rect 24952 12112 25004 12164
rect 30472 12180 30524 12232
rect 28264 12112 28316 12164
rect 31024 12112 31076 12164
rect 32220 12248 32272 12300
rect 32956 12316 33008 12368
rect 36636 12359 36688 12368
rect 32772 12291 32824 12300
rect 32772 12257 32781 12291
rect 32781 12257 32815 12291
rect 32815 12257 32824 12291
rect 32772 12248 32824 12257
rect 34336 12291 34388 12300
rect 34336 12257 34345 12291
rect 34345 12257 34379 12291
rect 34379 12257 34388 12291
rect 34336 12248 34388 12257
rect 36176 12291 36228 12300
rect 31208 12180 31260 12232
rect 32588 12180 32640 12232
rect 33784 12180 33836 12232
rect 33968 12180 34020 12232
rect 36176 12257 36185 12291
rect 36185 12257 36219 12291
rect 36219 12257 36228 12291
rect 36176 12248 36228 12257
rect 36636 12325 36645 12359
rect 36645 12325 36679 12359
rect 36679 12325 36688 12359
rect 36636 12316 36688 12325
rect 41144 12316 41196 12368
rect 44548 12359 44600 12368
rect 34980 12180 35032 12232
rect 36452 12180 36504 12232
rect 37832 12180 37884 12232
rect 38752 12223 38804 12232
rect 38752 12189 38761 12223
rect 38761 12189 38795 12223
rect 38795 12189 38804 12223
rect 38752 12180 38804 12189
rect 39028 12223 39080 12232
rect 39028 12189 39037 12223
rect 39037 12189 39071 12223
rect 39071 12189 39080 12223
rect 39028 12180 39080 12189
rect 41420 12248 41472 12300
rect 41512 12248 41564 12300
rect 42064 12291 42116 12300
rect 42064 12257 42073 12291
rect 42073 12257 42107 12291
rect 42107 12257 42116 12291
rect 42064 12248 42116 12257
rect 42248 12248 42300 12300
rect 44548 12325 44557 12359
rect 44557 12325 44591 12359
rect 44591 12325 44600 12359
rect 44548 12316 44600 12325
rect 47124 12359 47176 12368
rect 47124 12325 47133 12359
rect 47133 12325 47167 12359
rect 47167 12325 47176 12359
rect 47124 12316 47176 12325
rect 50528 12316 50580 12368
rect 45192 12291 45244 12300
rect 45192 12257 45201 12291
rect 45201 12257 45235 12291
rect 45235 12257 45244 12291
rect 45192 12248 45244 12257
rect 45560 12291 45612 12300
rect 45560 12257 45569 12291
rect 45569 12257 45603 12291
rect 45603 12257 45612 12291
rect 45560 12248 45612 12257
rect 45836 12248 45888 12300
rect 41972 12180 42024 12232
rect 42156 12223 42208 12232
rect 42156 12189 42165 12223
rect 42165 12189 42199 12223
rect 42199 12189 42208 12223
rect 42156 12180 42208 12189
rect 44732 12180 44784 12232
rect 46572 12223 46624 12232
rect 46572 12189 46581 12223
rect 46581 12189 46615 12223
rect 46615 12189 46624 12223
rect 46572 12180 46624 12189
rect 43444 12112 43496 12164
rect 43812 12112 43864 12164
rect 46204 12112 46256 12164
rect 48228 12248 48280 12300
rect 50896 12291 50948 12300
rect 50896 12257 50905 12291
rect 50905 12257 50939 12291
rect 50939 12257 50948 12291
rect 50896 12248 50948 12257
rect 52552 12316 52604 12368
rect 53196 12384 53248 12436
rect 55036 12384 55088 12436
rect 54576 12359 54628 12368
rect 54576 12325 54585 12359
rect 54585 12325 54619 12359
rect 54619 12325 54628 12359
rect 54576 12316 54628 12325
rect 53472 12291 53524 12300
rect 53472 12257 53481 12291
rect 53481 12257 53515 12291
rect 53515 12257 53524 12291
rect 53472 12248 53524 12257
rect 53564 12248 53616 12300
rect 55864 12316 55916 12368
rect 55036 12248 55088 12300
rect 55772 12291 55824 12300
rect 53748 12180 53800 12232
rect 55220 12112 55272 12164
rect 55772 12257 55781 12291
rect 55781 12257 55815 12291
rect 55815 12257 55824 12291
rect 55772 12248 55824 12257
rect 58164 12291 58216 12300
rect 58164 12257 58173 12291
rect 58173 12257 58207 12291
rect 58207 12257 58216 12291
rect 58164 12248 58216 12257
rect 56048 12180 56100 12232
rect 59728 12248 59780 12300
rect 59084 12180 59136 12232
rect 58440 12112 58492 12164
rect 7288 12044 7340 12096
rect 8208 12044 8260 12096
rect 12992 12044 13044 12096
rect 13360 12044 13412 12096
rect 13544 12044 13596 12096
rect 14004 12044 14056 12096
rect 15108 12044 15160 12096
rect 15384 12044 15436 12096
rect 23572 12044 23624 12096
rect 23664 12044 23716 12096
rect 25504 12087 25556 12096
rect 25504 12053 25513 12087
rect 25513 12053 25547 12087
rect 25547 12053 25556 12087
rect 25504 12044 25556 12053
rect 34244 12044 34296 12096
rect 34428 12044 34480 12096
rect 35900 12044 35952 12096
rect 36728 12044 36780 12096
rect 37188 12044 37240 12096
rect 39672 12044 39724 12096
rect 40132 12087 40184 12096
rect 40132 12053 40141 12087
rect 40141 12053 40175 12087
rect 40175 12053 40184 12087
rect 40132 12044 40184 12053
rect 40684 12044 40736 12096
rect 50252 12044 50304 12096
rect 56232 12044 56284 12096
rect 11163 11942 11215 11994
rect 11227 11942 11279 11994
rect 11291 11942 11343 11994
rect 11355 11942 11407 11994
rect 31526 11942 31578 11994
rect 31590 11942 31642 11994
rect 31654 11942 31706 11994
rect 31718 11942 31770 11994
rect 51888 11942 51940 11994
rect 51952 11942 52004 11994
rect 52016 11942 52068 11994
rect 52080 11942 52132 11994
rect 7196 11840 7248 11892
rect 13176 11840 13228 11892
rect 13268 11840 13320 11892
rect 19892 11840 19944 11892
rect 20076 11883 20128 11892
rect 20076 11849 20085 11883
rect 20085 11849 20119 11883
rect 20119 11849 20128 11883
rect 20076 11840 20128 11849
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 3148 11679 3200 11688
rect 3148 11645 3157 11679
rect 3157 11645 3191 11679
rect 3191 11645 3200 11679
rect 3148 11636 3200 11645
rect 5080 11679 5132 11688
rect 5080 11645 5089 11679
rect 5089 11645 5123 11679
rect 5123 11645 5132 11679
rect 5080 11636 5132 11645
rect 5448 11636 5500 11688
rect 6920 11636 6972 11688
rect 7564 11747 7616 11756
rect 7564 11713 7573 11747
rect 7573 11713 7607 11747
rect 7607 11713 7616 11747
rect 7564 11704 7616 11713
rect 12348 11772 12400 11824
rect 12716 11772 12768 11824
rect 14372 11772 14424 11824
rect 21548 11840 21600 11892
rect 22100 11840 22152 11892
rect 25504 11840 25556 11892
rect 7932 11747 7984 11756
rect 7932 11713 7941 11747
rect 7941 11713 7975 11747
rect 7975 11713 7984 11747
rect 7932 11704 7984 11713
rect 11244 11704 11296 11756
rect 11520 11747 11572 11756
rect 11520 11713 11529 11747
rect 11529 11713 11563 11747
rect 11563 11713 11572 11747
rect 11520 11704 11572 11713
rect 12440 11704 12492 11756
rect 13360 11704 13412 11756
rect 13636 11704 13688 11756
rect 8024 11636 8076 11688
rect 8208 11636 8260 11688
rect 9036 11679 9088 11688
rect 9036 11645 9045 11679
rect 9045 11645 9079 11679
rect 9079 11645 9088 11679
rect 9036 11636 9088 11645
rect 11060 11679 11112 11688
rect 11060 11645 11069 11679
rect 11069 11645 11103 11679
rect 11103 11645 11112 11679
rect 11060 11636 11112 11645
rect 11336 11636 11388 11688
rect 13268 11636 13320 11688
rect 15016 11704 15068 11756
rect 14924 11679 14976 11688
rect 14924 11645 14933 11679
rect 14933 11645 14967 11679
rect 14967 11645 14976 11679
rect 14924 11636 14976 11645
rect 15384 11747 15436 11756
rect 15384 11713 15393 11747
rect 15393 11713 15427 11747
rect 15427 11713 15436 11747
rect 15384 11704 15436 11713
rect 20260 11704 20312 11756
rect 16212 11636 16264 11688
rect 14464 11611 14516 11620
rect 14464 11577 14473 11611
rect 14473 11577 14507 11611
rect 14507 11577 14516 11611
rect 14464 11568 14516 11577
rect 14556 11568 14608 11620
rect 19708 11636 19760 11688
rect 23756 11772 23808 11824
rect 28356 11772 28408 11824
rect 30196 11772 30248 11824
rect 20812 11704 20864 11756
rect 21088 11747 21140 11756
rect 21088 11713 21097 11747
rect 21097 11713 21131 11747
rect 21131 11713 21140 11747
rect 21088 11704 21140 11713
rect 21732 11704 21784 11756
rect 17500 11568 17552 11620
rect 18788 11611 18840 11620
rect 18788 11577 18797 11611
rect 18797 11577 18831 11611
rect 18831 11577 18840 11611
rect 18788 11568 18840 11577
rect 19340 11568 19392 11620
rect 12808 11500 12860 11552
rect 15752 11500 15804 11552
rect 16304 11543 16356 11552
rect 16304 11509 16313 11543
rect 16313 11509 16347 11543
rect 16347 11509 16356 11543
rect 16304 11500 16356 11509
rect 20628 11500 20680 11552
rect 23480 11636 23532 11688
rect 27344 11704 27396 11756
rect 24032 11636 24084 11688
rect 24768 11679 24820 11688
rect 24768 11645 24777 11679
rect 24777 11645 24811 11679
rect 24811 11645 24820 11679
rect 24768 11636 24820 11645
rect 25780 11636 25832 11688
rect 26148 11636 26200 11688
rect 26792 11636 26844 11688
rect 27620 11704 27672 11756
rect 27896 11704 27948 11756
rect 28080 11747 28132 11756
rect 28080 11713 28089 11747
rect 28089 11713 28123 11747
rect 28123 11713 28132 11747
rect 28080 11704 28132 11713
rect 20904 11568 20956 11620
rect 22468 11500 22520 11552
rect 27344 11568 27396 11620
rect 27804 11636 27856 11688
rect 30196 11679 30248 11688
rect 29828 11568 29880 11620
rect 25320 11500 25372 11552
rect 26056 11500 26108 11552
rect 27988 11500 28040 11552
rect 30196 11645 30205 11679
rect 30205 11645 30239 11679
rect 30239 11645 30248 11679
rect 30196 11636 30248 11645
rect 30748 11704 30800 11756
rect 32404 11840 32456 11892
rect 34336 11840 34388 11892
rect 38936 11840 38988 11892
rect 40132 11840 40184 11892
rect 45192 11840 45244 11892
rect 49700 11840 49752 11892
rect 32220 11636 32272 11688
rect 32404 11679 32456 11688
rect 32404 11645 32413 11679
rect 32413 11645 32447 11679
rect 32447 11645 32456 11679
rect 32404 11636 32456 11645
rect 32588 11747 32640 11756
rect 32588 11713 32597 11747
rect 32597 11713 32631 11747
rect 32631 11713 32640 11747
rect 32588 11704 32640 11713
rect 33692 11704 33744 11756
rect 33968 11747 34020 11756
rect 33968 11713 33977 11747
rect 33977 11713 34011 11747
rect 34011 11713 34020 11747
rect 33968 11704 34020 11713
rect 37372 11772 37424 11824
rect 41604 11772 41656 11824
rect 43720 11772 43772 11824
rect 33508 11636 33560 11688
rect 34152 11636 34204 11688
rect 34796 11704 34848 11756
rect 41236 11704 41288 11756
rect 41420 11704 41472 11756
rect 41972 11704 42024 11756
rect 44364 11704 44416 11756
rect 45284 11772 45336 11824
rect 46664 11772 46716 11824
rect 49240 11772 49292 11824
rect 52000 11815 52052 11824
rect 52000 11781 52009 11815
rect 52009 11781 52043 11815
rect 52043 11781 52052 11815
rect 52000 11772 52052 11781
rect 52920 11840 52972 11892
rect 55864 11840 55916 11892
rect 46296 11704 46348 11756
rect 56048 11772 56100 11824
rect 35716 11636 35768 11688
rect 36452 11636 36504 11688
rect 36636 11679 36688 11688
rect 36636 11645 36645 11679
rect 36645 11645 36679 11679
rect 36679 11645 36688 11679
rect 36636 11636 36688 11645
rect 36728 11636 36780 11688
rect 37096 11636 37148 11688
rect 41144 11636 41196 11688
rect 42340 11636 42392 11688
rect 30656 11568 30708 11620
rect 32772 11568 32824 11620
rect 34796 11568 34848 11620
rect 30840 11500 30892 11552
rect 33968 11500 34020 11552
rect 41420 11568 41472 11620
rect 42616 11636 42668 11688
rect 46204 11679 46256 11688
rect 42892 11568 42944 11620
rect 37648 11500 37700 11552
rect 42248 11500 42300 11552
rect 43168 11543 43220 11552
rect 43168 11509 43177 11543
rect 43177 11509 43211 11543
rect 43211 11509 43220 11543
rect 43168 11500 43220 11509
rect 46204 11645 46213 11679
rect 46213 11645 46247 11679
rect 46247 11645 46256 11679
rect 46204 11636 46256 11645
rect 48780 11679 48832 11688
rect 48780 11645 48789 11679
rect 48789 11645 48823 11679
rect 48823 11645 48832 11679
rect 48780 11636 48832 11645
rect 45192 11568 45244 11620
rect 48688 11568 48740 11620
rect 49700 11636 49752 11688
rect 50528 11679 50580 11688
rect 50528 11645 50537 11679
rect 50537 11645 50571 11679
rect 50571 11645 50580 11679
rect 50528 11636 50580 11645
rect 51632 11636 51684 11688
rect 55312 11704 55364 11756
rect 60464 11840 60516 11892
rect 53196 11636 53248 11688
rect 56784 11704 56836 11756
rect 56232 11679 56284 11688
rect 50620 11568 50672 11620
rect 49976 11500 50028 11552
rect 50528 11500 50580 11552
rect 51080 11500 51132 11552
rect 52368 11500 52420 11552
rect 56232 11645 56241 11679
rect 56241 11645 56275 11679
rect 56275 11645 56284 11679
rect 56232 11636 56284 11645
rect 56600 11636 56652 11688
rect 57336 11636 57388 11688
rect 56692 11568 56744 11620
rect 54668 11500 54720 11552
rect 56232 11500 56284 11552
rect 21344 11398 21396 11450
rect 21408 11398 21460 11450
rect 21472 11398 21524 11450
rect 21536 11398 21588 11450
rect 41707 11398 41759 11450
rect 41771 11398 41823 11450
rect 41835 11398 41887 11450
rect 41899 11398 41951 11450
rect 5080 11296 5132 11348
rect 6920 11271 6972 11280
rect 6920 11237 6929 11271
rect 6929 11237 6963 11271
rect 6963 11237 6972 11271
rect 6920 11228 6972 11237
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2780 11160 2832 11169
rect 3976 11160 4028 11212
rect 11336 11271 11388 11280
rect 3056 11092 3108 11144
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 4436 11024 4488 11076
rect 5540 11024 5592 11076
rect 6828 11092 6880 11144
rect 9036 11160 9088 11212
rect 10784 11203 10836 11212
rect 10784 11169 10793 11203
rect 10793 11169 10827 11203
rect 10827 11169 10836 11203
rect 10784 11160 10836 11169
rect 7472 11024 7524 11076
rect 10968 11160 11020 11212
rect 11336 11237 11345 11271
rect 11345 11237 11379 11271
rect 11379 11237 11388 11271
rect 11336 11228 11388 11237
rect 13176 11296 13228 11348
rect 14372 11228 14424 11280
rect 14924 11228 14976 11280
rect 14004 11160 14056 11212
rect 14096 11160 14148 11212
rect 16028 11160 16080 11212
rect 12164 11135 12216 11144
rect 12164 11101 12173 11135
rect 12173 11101 12207 11135
rect 12207 11101 12216 11135
rect 12164 11092 12216 11101
rect 15108 11092 15160 11144
rect 15200 11092 15252 11144
rect 21088 11296 21140 11348
rect 21640 11296 21692 11348
rect 18236 11228 18288 11280
rect 18788 11228 18840 11280
rect 19340 11203 19392 11212
rect 13452 11024 13504 11076
rect 16120 11024 16172 11076
rect 19340 11169 19349 11203
rect 19349 11169 19383 11203
rect 19383 11169 19392 11203
rect 19340 11160 19392 11169
rect 19708 11203 19760 11212
rect 19708 11169 19717 11203
rect 19717 11169 19751 11203
rect 19751 11169 19760 11203
rect 19708 11160 19760 11169
rect 20628 11228 20680 11280
rect 19892 11160 19944 11212
rect 19248 11092 19300 11144
rect 19616 11092 19668 11144
rect 20260 11092 20312 11144
rect 20904 11135 20956 11144
rect 20904 11101 20913 11135
rect 20913 11101 20947 11135
rect 20947 11101 20956 11135
rect 20904 11092 20956 11101
rect 22652 11160 22704 11212
rect 23296 11203 23348 11212
rect 23296 11169 23305 11203
rect 23305 11169 23339 11203
rect 23339 11169 23348 11203
rect 23296 11160 23348 11169
rect 24216 11203 24268 11212
rect 24216 11169 24225 11203
rect 24225 11169 24259 11203
rect 24259 11169 24268 11203
rect 24216 11160 24268 11169
rect 29828 11339 29880 11348
rect 29828 11305 29837 11339
rect 29837 11305 29871 11339
rect 29871 11305 29880 11339
rect 29828 11296 29880 11305
rect 30932 11296 30984 11348
rect 31116 11339 31168 11348
rect 31116 11305 31125 11339
rect 31125 11305 31159 11339
rect 31159 11305 31168 11339
rect 31116 11296 31168 11305
rect 32312 11339 32364 11348
rect 32312 11305 32321 11339
rect 32321 11305 32355 11339
rect 32355 11305 32364 11339
rect 32312 11296 32364 11305
rect 27160 11228 27212 11280
rect 28264 11228 28316 11280
rect 26056 11160 26108 11212
rect 27620 11160 27672 11212
rect 27896 11160 27948 11212
rect 28356 11203 28408 11212
rect 28356 11169 28365 11203
rect 28365 11169 28399 11203
rect 28399 11169 28408 11203
rect 28356 11160 28408 11169
rect 27804 11092 27856 11144
rect 29000 11160 29052 11212
rect 30196 11160 30248 11212
rect 30472 11160 30524 11212
rect 34244 11228 34296 11280
rect 40500 11296 40552 11348
rect 41420 11296 41472 11348
rect 47492 11296 47544 11348
rect 33508 11135 33560 11144
rect 21732 11024 21784 11076
rect 29000 11024 29052 11076
rect 9680 10956 9732 11008
rect 10876 10956 10928 11008
rect 12440 10956 12492 11008
rect 17500 10956 17552 11008
rect 22560 10956 22612 11008
rect 23388 10999 23440 11008
rect 23388 10965 23397 10999
rect 23397 10965 23431 10999
rect 23431 10965 23440 10999
rect 23388 10956 23440 10965
rect 26700 10956 26752 11008
rect 27068 10999 27120 11008
rect 27068 10965 27077 10999
rect 27077 10965 27111 10999
rect 27111 10965 27120 10999
rect 27068 10956 27120 10965
rect 33508 11101 33517 11135
rect 33517 11101 33551 11135
rect 33551 11101 33560 11135
rect 33508 11092 33560 11101
rect 33968 11160 34020 11212
rect 35072 11160 35124 11212
rect 36268 11203 36320 11212
rect 36268 11169 36277 11203
rect 36277 11169 36311 11203
rect 36311 11169 36320 11203
rect 36268 11160 36320 11169
rect 36544 11160 36596 11212
rect 36820 11160 36872 11212
rect 41420 11160 41472 11212
rect 34980 11092 35032 11144
rect 36636 11024 36688 11076
rect 33600 10956 33652 11008
rect 34888 10956 34940 11008
rect 36452 10956 36504 11008
rect 38752 11092 38804 11144
rect 39212 11135 39264 11144
rect 39212 11101 39221 11135
rect 39221 11101 39255 11135
rect 39255 11101 39264 11135
rect 39212 11092 39264 11101
rect 39488 11135 39540 11144
rect 39488 11101 39497 11135
rect 39497 11101 39531 11135
rect 39531 11101 39540 11135
rect 39488 11092 39540 11101
rect 41328 11092 41380 11144
rect 42616 11160 42668 11212
rect 43168 11160 43220 11212
rect 43812 11160 43864 11212
rect 44088 11228 44140 11280
rect 48044 11271 48096 11280
rect 48044 11237 48053 11271
rect 48053 11237 48087 11271
rect 48087 11237 48096 11271
rect 48044 11228 48096 11237
rect 49056 11160 49108 11212
rect 49240 11203 49292 11212
rect 49240 11169 49249 11203
rect 49249 11169 49283 11203
rect 49283 11169 49292 11203
rect 49240 11160 49292 11169
rect 51540 11296 51592 11348
rect 50620 11271 50672 11280
rect 50620 11237 50629 11271
rect 50629 11237 50663 11271
rect 50663 11237 50672 11271
rect 50620 11228 50672 11237
rect 53196 11296 53248 11348
rect 53748 11228 53800 11280
rect 52000 11203 52052 11212
rect 44824 11092 44876 11144
rect 45192 11092 45244 11144
rect 46112 11092 46164 11144
rect 47492 11135 47544 11144
rect 47492 11101 47501 11135
rect 47501 11101 47535 11135
rect 47535 11101 47544 11135
rect 47492 11092 47544 11101
rect 51540 11092 51592 11144
rect 52000 11169 52009 11203
rect 52009 11169 52043 11203
rect 52043 11169 52052 11203
rect 52000 11160 52052 11169
rect 54668 11203 54720 11212
rect 54668 11169 54677 11203
rect 54677 11169 54711 11203
rect 54711 11169 54720 11203
rect 54668 11160 54720 11169
rect 56324 11296 56376 11348
rect 59084 11339 59136 11348
rect 59084 11305 59093 11339
rect 59093 11305 59127 11339
rect 59127 11305 59136 11339
rect 59084 11296 59136 11305
rect 56692 11203 56744 11212
rect 38844 11024 38896 11076
rect 54576 11135 54628 11144
rect 54576 11101 54585 11135
rect 54585 11101 54619 11135
rect 54619 11101 54628 11135
rect 54576 11092 54628 11101
rect 43536 10956 43588 11008
rect 43812 10956 43864 11008
rect 56232 11024 56284 11076
rect 46572 10956 46624 11008
rect 46940 10956 46992 11008
rect 48412 10956 48464 11008
rect 54576 10956 54628 11008
rect 56692 11169 56701 11203
rect 56701 11169 56735 11203
rect 56735 11169 56744 11203
rect 56692 11160 56744 11169
rect 56600 11092 56652 11144
rect 57336 10956 57388 11008
rect 11163 10854 11215 10906
rect 11227 10854 11279 10906
rect 11291 10854 11343 10906
rect 11355 10854 11407 10906
rect 31526 10854 31578 10906
rect 31590 10854 31642 10906
rect 31654 10854 31706 10906
rect 31718 10854 31770 10906
rect 51888 10854 51940 10906
rect 51952 10854 52004 10906
rect 52016 10854 52068 10906
rect 52080 10854 52132 10906
rect 3148 10752 3200 10804
rect 6644 10752 6696 10804
rect 7104 10795 7156 10804
rect 5448 10616 5500 10668
rect 7104 10761 7113 10795
rect 7113 10761 7147 10795
rect 7147 10761 7156 10795
rect 7104 10752 7156 10761
rect 7564 10752 7616 10804
rect 9680 10752 9732 10804
rect 18420 10752 18472 10804
rect 15016 10684 15068 10736
rect 16396 10727 16448 10736
rect 16396 10693 16405 10727
rect 16405 10693 16439 10727
rect 16439 10693 16448 10727
rect 16396 10684 16448 10693
rect 16672 10684 16724 10736
rect 2780 10548 2832 10600
rect 3976 10548 4028 10600
rect 6736 10548 6788 10600
rect 8760 10591 8812 10600
rect 8760 10557 8769 10591
rect 8769 10557 8803 10591
rect 8803 10557 8812 10591
rect 8760 10548 8812 10557
rect 9864 10591 9916 10600
rect 9864 10557 9873 10591
rect 9873 10557 9907 10591
rect 9907 10557 9916 10591
rect 9864 10548 9916 10557
rect 10968 10591 11020 10600
rect 10968 10557 10977 10591
rect 10977 10557 11011 10591
rect 11011 10557 11020 10591
rect 10968 10548 11020 10557
rect 12164 10616 12216 10668
rect 14464 10616 14516 10668
rect 20904 10752 20956 10804
rect 32312 10752 32364 10804
rect 20628 10684 20680 10736
rect 11612 10548 11664 10600
rect 15292 10591 15344 10600
rect 4068 10412 4120 10464
rect 12072 10480 12124 10532
rect 7288 10412 7340 10464
rect 7656 10412 7708 10464
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 10968 10412 11020 10464
rect 13176 10412 13228 10464
rect 15292 10557 15301 10591
rect 15301 10557 15335 10591
rect 15335 10557 15344 10591
rect 15292 10548 15344 10557
rect 16304 10548 16356 10600
rect 19340 10591 19392 10600
rect 19340 10557 19349 10591
rect 19349 10557 19383 10591
rect 19383 10557 19392 10591
rect 19616 10616 19668 10668
rect 19340 10548 19392 10557
rect 19708 10548 19760 10600
rect 22192 10616 22244 10668
rect 24216 10616 24268 10668
rect 24768 10616 24820 10668
rect 25872 10616 25924 10668
rect 27068 10616 27120 10668
rect 27620 10616 27672 10668
rect 20812 10591 20864 10600
rect 20812 10557 20821 10591
rect 20821 10557 20855 10591
rect 20855 10557 20864 10591
rect 20812 10548 20864 10557
rect 23572 10548 23624 10600
rect 19248 10523 19300 10532
rect 19248 10489 19257 10523
rect 19257 10489 19291 10523
rect 19291 10489 19300 10523
rect 19248 10480 19300 10489
rect 15752 10412 15804 10464
rect 16396 10412 16448 10464
rect 18972 10412 19024 10464
rect 19064 10412 19116 10464
rect 19432 10412 19484 10464
rect 20168 10412 20220 10464
rect 22560 10480 22612 10532
rect 23848 10455 23900 10464
rect 23848 10421 23857 10455
rect 23857 10421 23891 10455
rect 23891 10421 23900 10455
rect 23848 10412 23900 10421
rect 25412 10548 25464 10600
rect 30104 10548 30156 10600
rect 30656 10591 30708 10600
rect 30656 10557 30665 10591
rect 30665 10557 30699 10591
rect 30699 10557 30708 10591
rect 30656 10548 30708 10557
rect 31852 10591 31904 10600
rect 31852 10557 31861 10591
rect 31861 10557 31895 10591
rect 31895 10557 31904 10591
rect 31852 10548 31904 10557
rect 33140 10548 33192 10600
rect 33876 10684 33928 10736
rect 36084 10752 36136 10804
rect 43720 10795 43772 10804
rect 43720 10761 43729 10795
rect 43729 10761 43763 10795
rect 43763 10761 43772 10795
rect 43720 10752 43772 10761
rect 39028 10684 39080 10736
rect 39212 10616 39264 10668
rect 42340 10616 42392 10668
rect 45100 10659 45152 10668
rect 45100 10625 45109 10659
rect 45109 10625 45143 10659
rect 45143 10625 45152 10659
rect 45100 10616 45152 10625
rect 46112 10659 46164 10668
rect 46112 10625 46121 10659
rect 46121 10625 46155 10659
rect 46155 10625 46164 10659
rect 46112 10616 46164 10625
rect 49056 10752 49108 10804
rect 50068 10752 50120 10804
rect 53104 10752 53156 10804
rect 56784 10684 56836 10736
rect 52368 10616 52420 10668
rect 57336 10659 57388 10668
rect 33784 10591 33836 10600
rect 33784 10557 33803 10591
rect 33803 10557 33836 10591
rect 33784 10548 33836 10557
rect 34888 10591 34940 10600
rect 34888 10557 34897 10591
rect 34897 10557 34931 10591
rect 34931 10557 34940 10591
rect 34888 10548 34940 10557
rect 38660 10591 38712 10600
rect 38660 10557 38669 10591
rect 38669 10557 38703 10591
rect 38703 10557 38712 10591
rect 38660 10548 38712 10557
rect 38844 10591 38896 10600
rect 38844 10557 38853 10591
rect 38853 10557 38887 10591
rect 38887 10557 38896 10591
rect 38844 10548 38896 10557
rect 38936 10548 38988 10600
rect 42432 10591 42484 10600
rect 42432 10557 42441 10591
rect 42441 10557 42475 10591
rect 42475 10557 42484 10591
rect 42432 10548 42484 10557
rect 44824 10591 44876 10600
rect 44824 10557 44833 10591
rect 44833 10557 44867 10591
rect 44867 10557 44876 10591
rect 44824 10548 44876 10557
rect 45928 10548 45980 10600
rect 46940 10591 46992 10600
rect 46940 10557 46949 10591
rect 46949 10557 46983 10591
rect 46983 10557 46992 10591
rect 46940 10548 46992 10557
rect 47216 10548 47268 10600
rect 48964 10548 49016 10600
rect 25780 10523 25832 10532
rect 25780 10489 25789 10523
rect 25789 10489 25823 10523
rect 25823 10489 25832 10523
rect 25780 10480 25832 10489
rect 27620 10480 27672 10532
rect 30472 10480 30524 10532
rect 48412 10480 48464 10532
rect 26148 10412 26200 10464
rect 26884 10412 26936 10464
rect 27528 10412 27580 10464
rect 30840 10455 30892 10464
rect 30840 10421 30849 10455
rect 30849 10421 30883 10455
rect 30883 10421 30892 10455
rect 30840 10412 30892 10421
rect 32036 10455 32088 10464
rect 32036 10421 32045 10455
rect 32045 10421 32079 10455
rect 32079 10421 32088 10455
rect 32036 10412 32088 10421
rect 46388 10412 46440 10464
rect 52920 10591 52972 10600
rect 49332 10480 49384 10532
rect 51356 10480 51408 10532
rect 52920 10557 52929 10591
rect 52929 10557 52963 10591
rect 52963 10557 52972 10591
rect 52920 10548 52972 10557
rect 57336 10625 57345 10659
rect 57345 10625 57379 10659
rect 57379 10625 57388 10659
rect 57336 10616 57388 10625
rect 54300 10591 54352 10600
rect 54300 10557 54309 10591
rect 54309 10557 54343 10591
rect 54343 10557 54352 10591
rect 54300 10548 54352 10557
rect 55404 10548 55456 10600
rect 56048 10591 56100 10600
rect 56048 10557 56057 10591
rect 56057 10557 56091 10591
rect 56091 10557 56100 10591
rect 56048 10548 56100 10557
rect 56232 10591 56284 10600
rect 56232 10557 56241 10591
rect 56241 10557 56275 10591
rect 56275 10557 56284 10591
rect 56232 10548 56284 10557
rect 53196 10480 53248 10532
rect 55772 10480 55824 10532
rect 51448 10412 51500 10464
rect 54760 10412 54812 10464
rect 58716 10455 58768 10464
rect 58716 10421 58725 10455
rect 58725 10421 58759 10455
rect 58759 10421 58768 10455
rect 58716 10412 58768 10421
rect 21344 10310 21396 10362
rect 21408 10310 21460 10362
rect 21472 10310 21524 10362
rect 21536 10310 21588 10362
rect 41707 10310 41759 10362
rect 41771 10310 41823 10362
rect 41835 10310 41887 10362
rect 41899 10310 41951 10362
rect 5080 10208 5132 10260
rect 10784 10208 10836 10260
rect 11796 10208 11848 10260
rect 12256 10208 12308 10260
rect 7012 10140 7064 10192
rect 13728 10140 13780 10192
rect 15108 10140 15160 10192
rect 15384 10140 15436 10192
rect 19248 10208 19300 10260
rect 29736 10208 29788 10260
rect 34980 10251 35032 10260
rect 34980 10217 34989 10251
rect 34989 10217 35023 10251
rect 35023 10217 35032 10251
rect 34980 10208 35032 10217
rect 36360 10251 36412 10260
rect 36360 10217 36369 10251
rect 36369 10217 36403 10251
rect 36403 10217 36412 10251
rect 36360 10208 36412 10217
rect 19616 10183 19668 10192
rect 19616 10149 19625 10183
rect 19625 10149 19659 10183
rect 19659 10149 19668 10183
rect 19616 10140 19668 10149
rect 24768 10140 24820 10192
rect 6644 10115 6696 10124
rect 6644 10081 6653 10115
rect 6653 10081 6687 10115
rect 6687 10081 6696 10115
rect 6644 10072 6696 10081
rect 10048 10115 10100 10124
rect 10048 10081 10057 10115
rect 10057 10081 10091 10115
rect 10091 10081 10100 10115
rect 10048 10072 10100 10081
rect 11612 10072 11664 10124
rect 11888 10072 11940 10124
rect 12072 10115 12124 10124
rect 12072 10081 12081 10115
rect 12081 10081 12115 10115
rect 12115 10081 12124 10115
rect 12072 10072 12124 10081
rect 3976 10004 4028 10056
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 9680 10004 9732 10056
rect 10876 10004 10928 10056
rect 13360 10072 13412 10124
rect 13176 10004 13228 10056
rect 15016 10072 15068 10124
rect 15844 10072 15896 10124
rect 16120 10115 16172 10124
rect 16120 10081 16129 10115
rect 16129 10081 16163 10115
rect 16163 10081 16172 10115
rect 16120 10072 16172 10081
rect 18420 10072 18472 10124
rect 19432 10115 19484 10124
rect 19432 10081 19441 10115
rect 19441 10081 19475 10115
rect 19475 10081 19484 10115
rect 19432 10072 19484 10081
rect 21088 10115 21140 10124
rect 21088 10081 21097 10115
rect 21097 10081 21131 10115
rect 21131 10081 21140 10115
rect 21088 10072 21140 10081
rect 21272 10072 21324 10124
rect 21824 10072 21876 10124
rect 13820 10047 13872 10056
rect 13820 10013 13829 10047
rect 13829 10013 13863 10047
rect 13863 10013 13872 10047
rect 13820 10004 13872 10013
rect 17592 10004 17644 10056
rect 19340 10004 19392 10056
rect 22192 10115 22244 10124
rect 22192 10081 22201 10115
rect 22201 10081 22235 10115
rect 22235 10081 22244 10115
rect 22192 10072 22244 10081
rect 23388 10072 23440 10124
rect 23572 10072 23624 10124
rect 25780 10140 25832 10192
rect 39488 10140 39540 10192
rect 41420 10140 41472 10192
rect 25044 10115 25096 10124
rect 25044 10081 25053 10115
rect 25053 10081 25087 10115
rect 25087 10081 25096 10115
rect 25044 10072 25096 10081
rect 26424 10072 26476 10124
rect 26884 10072 26936 10124
rect 27068 10115 27120 10124
rect 27068 10081 27077 10115
rect 27077 10081 27111 10115
rect 27111 10081 27120 10115
rect 27068 10072 27120 10081
rect 27620 10072 27672 10124
rect 29000 10115 29052 10124
rect 11704 9936 11756 9988
rect 12072 9936 12124 9988
rect 13452 9936 13504 9988
rect 19616 9936 19668 9988
rect 21272 9979 21324 9988
rect 21272 9945 21281 9979
rect 21281 9945 21315 9979
rect 21315 9945 21324 9979
rect 21272 9936 21324 9945
rect 10232 9911 10284 9920
rect 10232 9877 10241 9911
rect 10241 9877 10275 9911
rect 10275 9877 10284 9911
rect 10232 9868 10284 9877
rect 11520 9868 11572 9920
rect 13728 9911 13780 9920
rect 13728 9877 13737 9911
rect 13737 9877 13771 9911
rect 13771 9877 13780 9911
rect 13728 9868 13780 9877
rect 16028 9868 16080 9920
rect 21180 9868 21232 9920
rect 24676 10004 24728 10056
rect 25320 10004 25372 10056
rect 29000 10081 29009 10115
rect 29009 10081 29043 10115
rect 29043 10081 29052 10115
rect 29000 10072 29052 10081
rect 30656 10072 30708 10124
rect 32128 10072 32180 10124
rect 32312 10115 32364 10124
rect 32312 10081 32321 10115
rect 32321 10081 32355 10115
rect 32355 10081 32364 10115
rect 32312 10072 32364 10081
rect 33600 10115 33652 10124
rect 33600 10081 33609 10115
rect 33609 10081 33643 10115
rect 33643 10081 33652 10115
rect 33600 10072 33652 10081
rect 34152 10072 34204 10124
rect 37740 10115 37792 10124
rect 37740 10081 37749 10115
rect 37749 10081 37783 10115
rect 37783 10081 37792 10115
rect 37740 10072 37792 10081
rect 39580 10072 39632 10124
rect 32220 10047 32272 10056
rect 32220 10013 32229 10047
rect 32229 10013 32263 10047
rect 32263 10013 32272 10047
rect 32220 10004 32272 10013
rect 33416 10004 33468 10056
rect 35624 10004 35676 10056
rect 38844 10004 38896 10056
rect 40500 10072 40552 10124
rect 41604 10072 41656 10124
rect 43720 10140 43772 10192
rect 42156 10115 42208 10124
rect 42156 10081 42165 10115
rect 42165 10081 42199 10115
rect 42199 10081 42208 10115
rect 42156 10072 42208 10081
rect 23296 9936 23348 9988
rect 26700 9936 26752 9988
rect 27436 9936 27488 9988
rect 27712 9936 27764 9988
rect 42432 9936 42484 9988
rect 22928 9868 22980 9920
rect 25044 9868 25096 9920
rect 27620 9868 27672 9920
rect 36912 9868 36964 9920
rect 44916 10208 44968 10260
rect 47492 10208 47544 10260
rect 47216 10140 47268 10192
rect 49332 10208 49384 10260
rect 48964 10183 49016 10192
rect 48964 10149 48973 10183
rect 48973 10149 49007 10183
rect 49007 10149 49016 10183
rect 48964 10140 49016 10149
rect 55772 10183 55824 10192
rect 55772 10149 55781 10183
rect 55781 10149 55815 10183
rect 55815 10149 55824 10183
rect 55772 10140 55824 10149
rect 45100 10072 45152 10124
rect 46112 10072 46164 10124
rect 49516 10072 49568 10124
rect 50068 10072 50120 10124
rect 51356 10072 51408 10124
rect 54668 10115 54720 10124
rect 44640 10047 44692 10056
rect 44640 10013 44649 10047
rect 44649 10013 44683 10047
rect 44683 10013 44692 10047
rect 44640 10004 44692 10013
rect 49700 10004 49752 10056
rect 51540 10047 51592 10056
rect 51540 10013 51549 10047
rect 51549 10013 51583 10047
rect 51583 10013 51592 10047
rect 51540 10004 51592 10013
rect 51724 10004 51776 10056
rect 54668 10081 54677 10115
rect 54677 10081 54711 10115
rect 54711 10081 54720 10115
rect 54668 10072 54720 10081
rect 59360 10208 59412 10260
rect 54576 10004 54628 10056
rect 58716 10072 58768 10124
rect 56600 9936 56652 9988
rect 57336 10004 57388 10056
rect 58072 10004 58124 10056
rect 50252 9868 50304 9920
rect 53196 9868 53248 9920
rect 54852 9911 54904 9920
rect 54852 9877 54861 9911
rect 54861 9877 54895 9911
rect 54895 9877 54904 9911
rect 54852 9868 54904 9877
rect 58532 9868 58584 9920
rect 11163 9766 11215 9818
rect 11227 9766 11279 9818
rect 11291 9766 11343 9818
rect 11355 9766 11407 9818
rect 31526 9766 31578 9818
rect 31590 9766 31642 9818
rect 31654 9766 31706 9818
rect 31718 9766 31770 9818
rect 51888 9766 51940 9818
rect 51952 9766 52004 9818
rect 52016 9766 52068 9818
rect 52080 9766 52132 9818
rect 9864 9664 9916 9716
rect 13452 9664 13504 9716
rect 6736 9596 6788 9648
rect 15292 9596 15344 9648
rect 17500 9596 17552 9648
rect 3976 9528 4028 9580
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 2964 9324 3016 9376
rect 10968 9528 11020 9580
rect 12164 9528 12216 9580
rect 15844 9571 15896 9580
rect 15844 9537 15853 9571
rect 15853 9537 15887 9571
rect 15887 9537 15896 9571
rect 15844 9528 15896 9537
rect 7196 9460 7248 9512
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 7656 9503 7708 9512
rect 7656 9469 7665 9503
rect 7665 9469 7699 9503
rect 7699 9469 7708 9503
rect 7656 9460 7708 9469
rect 11060 9460 11112 9512
rect 11520 9460 11572 9512
rect 12716 9503 12768 9512
rect 12716 9469 12725 9503
rect 12725 9469 12759 9503
rect 12759 9469 12768 9503
rect 12716 9460 12768 9469
rect 12992 9460 13044 9512
rect 13728 9460 13780 9512
rect 15384 9503 15436 9512
rect 8668 9324 8720 9376
rect 13820 9392 13872 9444
rect 14648 9392 14700 9444
rect 15384 9469 15393 9503
rect 15393 9469 15427 9503
rect 15427 9469 15436 9503
rect 15384 9460 15436 9469
rect 16672 9528 16724 9580
rect 16580 9460 16632 9512
rect 19616 9596 19668 9648
rect 20720 9596 20772 9648
rect 23112 9596 23164 9648
rect 23756 9639 23808 9648
rect 23756 9605 23765 9639
rect 23765 9605 23799 9639
rect 23799 9605 23808 9639
rect 23756 9596 23808 9605
rect 24124 9596 24176 9648
rect 27896 9596 27948 9648
rect 33508 9596 33560 9648
rect 36268 9596 36320 9648
rect 44364 9664 44416 9716
rect 44916 9664 44968 9716
rect 45192 9664 45244 9716
rect 48136 9664 48188 9716
rect 48596 9664 48648 9716
rect 49056 9707 49108 9716
rect 49056 9673 49065 9707
rect 49065 9673 49099 9707
rect 49099 9673 49108 9707
rect 49056 9664 49108 9673
rect 37096 9596 37148 9648
rect 19524 9528 19576 9580
rect 18328 9503 18380 9512
rect 18328 9469 18337 9503
rect 18337 9469 18371 9503
rect 18371 9469 18380 9503
rect 18328 9460 18380 9469
rect 18420 9503 18472 9512
rect 18420 9469 18429 9503
rect 18429 9469 18463 9503
rect 18463 9469 18472 9503
rect 18420 9460 18472 9469
rect 19708 9503 19760 9512
rect 19708 9469 19717 9503
rect 19717 9469 19751 9503
rect 19751 9469 19760 9503
rect 19708 9460 19760 9469
rect 20904 9460 20956 9512
rect 21732 9460 21784 9512
rect 22192 9503 22244 9512
rect 22192 9469 22201 9503
rect 22201 9469 22235 9503
rect 22235 9469 22244 9503
rect 22192 9460 22244 9469
rect 23940 9528 23992 9580
rect 23204 9460 23256 9512
rect 24216 9460 24268 9512
rect 25320 9503 25372 9512
rect 25320 9469 25329 9503
rect 25329 9469 25363 9503
rect 25363 9469 25372 9503
rect 25320 9460 25372 9469
rect 26148 9528 26200 9580
rect 26424 9528 26476 9580
rect 27160 9528 27212 9580
rect 29736 9571 29788 9580
rect 27252 9503 27304 9512
rect 27252 9469 27261 9503
rect 27261 9469 27295 9503
rect 27295 9469 27304 9503
rect 27252 9460 27304 9469
rect 27528 9460 27580 9512
rect 9680 9324 9732 9376
rect 11796 9324 11848 9376
rect 18328 9324 18380 9376
rect 19340 9324 19392 9376
rect 21088 9392 21140 9444
rect 22008 9392 22060 9444
rect 26516 9392 26568 9444
rect 27068 9392 27120 9444
rect 29000 9460 29052 9512
rect 29736 9537 29745 9571
rect 29745 9537 29779 9571
rect 29779 9537 29788 9571
rect 29736 9528 29788 9537
rect 32404 9528 32456 9580
rect 37280 9528 37332 9580
rect 41512 9528 41564 9580
rect 42800 9596 42852 9648
rect 48504 9596 48556 9648
rect 48688 9596 48740 9648
rect 43260 9528 43312 9580
rect 43904 9528 43956 9580
rect 45560 9528 45612 9580
rect 46112 9571 46164 9580
rect 46112 9537 46121 9571
rect 46121 9537 46155 9571
rect 46155 9537 46164 9571
rect 46112 9528 46164 9537
rect 29276 9435 29328 9444
rect 29276 9401 29285 9435
rect 29285 9401 29319 9435
rect 29319 9401 29328 9435
rect 29276 9392 29328 9401
rect 30748 9435 30800 9444
rect 30748 9401 30757 9435
rect 30757 9401 30791 9435
rect 30791 9401 30800 9435
rect 30748 9392 30800 9401
rect 31852 9460 31904 9512
rect 32680 9460 32732 9512
rect 33416 9503 33468 9512
rect 33416 9469 33425 9503
rect 33425 9469 33459 9503
rect 33459 9469 33468 9503
rect 33416 9460 33468 9469
rect 33876 9503 33928 9512
rect 33876 9469 33885 9503
rect 33885 9469 33919 9503
rect 33919 9469 33928 9503
rect 35348 9503 35400 9512
rect 33876 9460 33928 9469
rect 20996 9324 21048 9376
rect 21640 9324 21692 9376
rect 27804 9324 27856 9376
rect 31300 9324 31352 9376
rect 32404 9324 32456 9376
rect 32772 9367 32824 9376
rect 32772 9333 32781 9367
rect 32781 9333 32815 9367
rect 32815 9333 32824 9367
rect 32772 9324 32824 9333
rect 33968 9392 34020 9444
rect 34980 9392 35032 9444
rect 34796 9324 34848 9376
rect 35348 9469 35357 9503
rect 35357 9469 35391 9503
rect 35391 9469 35400 9503
rect 35348 9460 35400 9469
rect 35440 9460 35492 9512
rect 35900 9460 35952 9512
rect 36452 9460 36504 9512
rect 36728 9503 36780 9512
rect 36728 9469 36737 9503
rect 36737 9469 36771 9503
rect 36771 9469 36780 9503
rect 36728 9460 36780 9469
rect 36636 9392 36688 9444
rect 38752 9460 38804 9512
rect 41420 9503 41472 9512
rect 37280 9392 37332 9444
rect 36820 9324 36872 9376
rect 41420 9469 41429 9503
rect 41429 9469 41463 9503
rect 41463 9469 41472 9503
rect 41420 9460 41472 9469
rect 41880 9460 41932 9512
rect 42064 9503 42116 9512
rect 42064 9469 42073 9503
rect 42073 9469 42107 9503
rect 42107 9469 42116 9503
rect 42064 9460 42116 9469
rect 44364 9460 44416 9512
rect 46388 9503 46440 9512
rect 46388 9469 46397 9503
rect 46397 9469 46431 9503
rect 46431 9469 46440 9503
rect 46388 9460 46440 9469
rect 47492 9460 47544 9512
rect 47768 9503 47820 9512
rect 47768 9469 47777 9503
rect 47777 9469 47811 9503
rect 47811 9469 47820 9503
rect 49240 9503 49292 9512
rect 47768 9460 47820 9469
rect 49240 9469 49249 9503
rect 49249 9469 49283 9503
rect 49283 9469 49292 9503
rect 49240 9460 49292 9469
rect 49792 9460 49844 9512
rect 50436 9503 50488 9512
rect 50436 9469 50445 9503
rect 50445 9469 50479 9503
rect 50479 9469 50488 9503
rect 50436 9460 50488 9469
rect 39304 9392 39356 9444
rect 39948 9324 40000 9376
rect 44088 9392 44140 9444
rect 46112 9392 46164 9444
rect 46480 9435 46532 9444
rect 46480 9401 46489 9435
rect 46489 9401 46523 9435
rect 46523 9401 46532 9435
rect 46848 9435 46900 9444
rect 46480 9392 46532 9401
rect 46848 9401 46857 9435
rect 46857 9401 46891 9435
rect 46891 9401 46900 9435
rect 46848 9392 46900 9401
rect 54852 9596 54904 9648
rect 54668 9528 54720 9580
rect 51264 9460 51316 9512
rect 51540 9460 51592 9512
rect 52736 9460 52788 9512
rect 54852 9460 54904 9512
rect 51724 9392 51776 9444
rect 54760 9392 54812 9444
rect 43352 9324 43404 9376
rect 45008 9324 45060 9376
rect 46204 9324 46256 9376
rect 49424 9324 49476 9376
rect 52920 9324 52972 9376
rect 54300 9324 54352 9376
rect 57336 9460 57388 9512
rect 57980 9460 58032 9512
rect 58348 9503 58400 9512
rect 58348 9469 58357 9503
rect 58357 9469 58391 9503
rect 58391 9469 58400 9503
rect 58348 9460 58400 9469
rect 55772 9435 55824 9444
rect 55772 9401 55781 9435
rect 55781 9401 55815 9435
rect 55815 9401 55824 9435
rect 55772 9392 55824 9401
rect 60188 9324 60240 9376
rect 21344 9222 21396 9274
rect 21408 9222 21460 9274
rect 21472 9222 21524 9274
rect 21536 9222 21588 9274
rect 41707 9222 41759 9274
rect 41771 9222 41823 9274
rect 41835 9222 41887 9274
rect 41899 9222 41951 9274
rect 388 9120 440 9172
rect 30748 9120 30800 9172
rect 32312 9120 32364 9172
rect 36636 9120 36688 9172
rect 36728 9120 36780 9172
rect 3240 9052 3292 9104
rect 4712 9095 4764 9104
rect 4712 9061 4721 9095
rect 4721 9061 4755 9095
rect 4755 9061 4764 9095
rect 4712 9052 4764 9061
rect 2872 8984 2924 9036
rect 2964 9027 3016 9036
rect 2964 8993 2973 9027
rect 2973 8993 3007 9027
rect 3007 8993 3016 9027
rect 2964 8984 3016 8993
rect 4528 8984 4580 9036
rect 5540 9027 5592 9036
rect 5540 8993 5549 9027
rect 5549 8993 5583 9027
rect 5583 8993 5592 9027
rect 5540 8984 5592 8993
rect 5632 9027 5684 9036
rect 5632 8993 5641 9027
rect 5641 8993 5675 9027
rect 5675 8993 5684 9027
rect 5632 8984 5684 8993
rect 7472 8984 7524 9036
rect 9588 9052 9640 9104
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 10600 8984 10652 9036
rect 11796 9052 11848 9104
rect 12348 9027 12400 9036
rect 12348 8993 12357 9027
rect 12357 8993 12391 9027
rect 12391 8993 12400 9027
rect 12348 8984 12400 8993
rect 13728 9027 13780 9036
rect 10784 8959 10836 8968
rect 10784 8925 10793 8959
rect 10793 8925 10827 8959
rect 10827 8925 10836 8959
rect 10784 8916 10836 8925
rect 11060 8916 11112 8968
rect 12256 8959 12308 8968
rect 12256 8925 12265 8959
rect 12265 8925 12299 8959
rect 12299 8925 12308 8959
rect 12256 8916 12308 8925
rect 8392 8780 8444 8832
rect 13728 8993 13737 9027
rect 13737 8993 13771 9027
rect 13771 8993 13780 9027
rect 13728 8984 13780 8993
rect 14280 9052 14332 9104
rect 17040 9095 17092 9104
rect 16396 8984 16448 9036
rect 17040 9061 17049 9095
rect 17049 9061 17083 9095
rect 17083 9061 17092 9095
rect 17040 9052 17092 9061
rect 18696 9052 18748 9104
rect 16488 8959 16540 8968
rect 16488 8925 16497 8959
rect 16497 8925 16531 8959
rect 16531 8925 16540 8959
rect 16488 8916 16540 8925
rect 18512 8984 18564 9036
rect 20720 9052 20772 9104
rect 20904 9095 20956 9104
rect 20904 9061 20913 9095
rect 20913 9061 20947 9095
rect 20947 9061 20956 9095
rect 20904 9052 20956 9061
rect 21824 9052 21876 9104
rect 24952 9052 25004 9104
rect 13820 8780 13872 8832
rect 15936 8780 15988 8832
rect 16120 8780 16172 8832
rect 17776 8916 17828 8968
rect 19616 8959 19668 8968
rect 19616 8925 19625 8959
rect 19625 8925 19659 8959
rect 19659 8925 19668 8959
rect 19616 8916 19668 8925
rect 20076 8916 20128 8968
rect 21180 8916 21232 8968
rect 21548 9027 21600 9036
rect 21548 8993 21557 9027
rect 21557 8993 21591 9027
rect 21591 8993 21600 9027
rect 21548 8984 21600 8993
rect 22284 8984 22336 9036
rect 23112 9027 23164 9036
rect 23112 8993 23121 9027
rect 23121 8993 23155 9027
rect 23155 8993 23164 9027
rect 23112 8984 23164 8993
rect 24768 9027 24820 9036
rect 21824 8916 21876 8968
rect 22100 8916 22152 8968
rect 24768 8993 24777 9027
rect 24777 8993 24811 9027
rect 24811 8993 24820 9027
rect 24768 8984 24820 8993
rect 27804 8984 27856 9036
rect 28908 9052 28960 9104
rect 35624 9095 35676 9104
rect 35624 9061 35633 9095
rect 35633 9061 35667 9095
rect 35667 9061 35676 9095
rect 35624 9052 35676 9061
rect 29184 8984 29236 9036
rect 30656 9027 30708 9036
rect 30656 8993 30665 9027
rect 30665 8993 30699 9027
rect 30699 8993 30708 9027
rect 30656 8984 30708 8993
rect 32128 9027 32180 9036
rect 32128 8993 32137 9027
rect 32137 8993 32171 9027
rect 32171 8993 32180 9027
rect 32128 8984 32180 8993
rect 32496 8984 32548 9036
rect 34888 8984 34940 9036
rect 37096 9052 37148 9104
rect 38660 9052 38712 9104
rect 36084 9027 36136 9036
rect 36084 8993 36093 9027
rect 36093 8993 36127 9027
rect 36127 8993 36136 9027
rect 36084 8984 36136 8993
rect 23664 8959 23716 8968
rect 17960 8848 18012 8900
rect 22376 8848 22428 8900
rect 22560 8848 22612 8900
rect 22744 8848 22796 8900
rect 23664 8925 23673 8959
rect 23673 8925 23707 8959
rect 23707 8925 23716 8959
rect 23664 8916 23716 8925
rect 24952 8916 25004 8968
rect 27344 8959 27396 8968
rect 27344 8925 27353 8959
rect 27353 8925 27387 8959
rect 27387 8925 27396 8959
rect 27344 8916 27396 8925
rect 27436 8916 27488 8968
rect 31300 8916 31352 8968
rect 32956 8916 33008 8968
rect 33416 8959 33468 8968
rect 33416 8925 33425 8959
rect 33425 8925 33459 8959
rect 33459 8925 33468 8959
rect 33416 8916 33468 8925
rect 35072 8916 35124 8968
rect 36820 8984 36872 9036
rect 39304 8984 39356 9036
rect 36728 8916 36780 8968
rect 23204 8848 23256 8900
rect 23848 8848 23900 8900
rect 19800 8780 19852 8832
rect 20812 8780 20864 8832
rect 20904 8780 20956 8832
rect 23388 8780 23440 8832
rect 25412 8780 25464 8832
rect 26608 8780 26660 8832
rect 29736 8780 29788 8832
rect 30196 8823 30248 8832
rect 30196 8789 30205 8823
rect 30205 8789 30239 8823
rect 30239 8789 30248 8823
rect 30196 8780 30248 8789
rect 30564 8780 30616 8832
rect 33048 8780 33100 8832
rect 37004 8848 37056 8900
rect 34796 8780 34848 8832
rect 37924 8848 37976 8900
rect 39948 8984 40000 9036
rect 41604 9052 41656 9104
rect 43260 9052 43312 9104
rect 43996 8959 44048 8968
rect 43996 8925 44005 8959
rect 44005 8925 44039 8959
rect 44039 8925 44048 8959
rect 43996 8916 44048 8925
rect 44272 8984 44324 9036
rect 44916 9027 44968 9036
rect 44916 8993 44925 9027
rect 44925 8993 44959 9027
rect 44959 8993 44968 9027
rect 44916 8984 44968 8993
rect 45652 9052 45704 9104
rect 45468 8984 45520 9036
rect 41328 8848 41380 8900
rect 45744 8916 45796 8968
rect 46940 8959 46992 8968
rect 46940 8925 46949 8959
rect 46949 8925 46983 8959
rect 46983 8925 46992 8959
rect 46940 8916 46992 8925
rect 47952 9027 48004 9036
rect 47952 8993 47961 9027
rect 47961 8993 47995 9027
rect 47995 8993 48004 9027
rect 47952 8984 48004 8993
rect 48688 8916 48740 8968
rect 49608 9027 49660 9036
rect 49608 8993 49617 9027
rect 49617 8993 49651 9027
rect 49651 8993 49660 9027
rect 49608 8984 49660 8993
rect 50436 8984 50488 9036
rect 51448 9027 51500 9036
rect 51448 8993 51457 9027
rect 51457 8993 51491 9027
rect 51491 8993 51500 9027
rect 51448 8984 51500 8993
rect 51724 8984 51776 9036
rect 52920 9052 52972 9104
rect 51356 8959 51408 8968
rect 37740 8780 37792 8832
rect 40040 8780 40092 8832
rect 44456 8780 44508 8832
rect 44824 8848 44876 8900
rect 47860 8848 47912 8900
rect 49608 8848 49660 8900
rect 51356 8925 51365 8959
rect 51365 8925 51399 8959
rect 51399 8925 51408 8959
rect 51356 8916 51408 8925
rect 54668 9052 54720 9104
rect 58348 9120 58400 9172
rect 58072 9095 58124 9104
rect 58072 9061 58081 9095
rect 58081 9061 58115 9095
rect 58115 9061 58124 9095
rect 58072 9052 58124 9061
rect 53656 8984 53708 9036
rect 54760 9027 54812 9036
rect 54760 8993 54769 9027
rect 54769 8993 54803 9027
rect 54803 8993 54812 9027
rect 54760 8984 54812 8993
rect 54944 8984 54996 9036
rect 56692 9027 56744 9036
rect 56692 8993 56701 9027
rect 56701 8993 56735 9027
rect 56735 8993 56744 9027
rect 56692 8984 56744 8993
rect 57060 9027 57112 9036
rect 57060 8993 57069 9027
rect 57069 8993 57103 9027
rect 57103 8993 57112 9027
rect 57060 8984 57112 8993
rect 57244 9027 57296 9036
rect 57244 8993 57253 9027
rect 57253 8993 57287 9027
rect 57287 8993 57296 9027
rect 57244 8984 57296 8993
rect 58716 9027 58768 9036
rect 53196 8959 53248 8968
rect 53196 8925 53205 8959
rect 53205 8925 53239 8959
rect 53239 8925 53248 8959
rect 53196 8916 53248 8925
rect 54852 8916 54904 8968
rect 58716 8993 58725 9027
rect 58725 8993 58759 9027
rect 58759 8993 58768 9027
rect 58716 8984 58768 8993
rect 59268 8984 59320 9036
rect 60188 9027 60240 9036
rect 60188 8993 60197 9027
rect 60197 8993 60231 9027
rect 60231 8993 60240 9027
rect 60188 8984 60240 8993
rect 58808 8959 58860 8968
rect 52184 8848 52236 8900
rect 45192 8780 45244 8832
rect 45836 8780 45888 8832
rect 49240 8780 49292 8832
rect 49424 8780 49476 8832
rect 55036 8848 55088 8900
rect 55312 8780 55364 8832
rect 58808 8925 58817 8959
rect 58817 8925 58851 8959
rect 58851 8925 58860 8959
rect 58808 8916 58860 8925
rect 59176 8959 59228 8968
rect 59176 8925 59185 8959
rect 59185 8925 59219 8959
rect 59219 8925 59228 8959
rect 59176 8916 59228 8925
rect 56876 8848 56928 8900
rect 11163 8678 11215 8730
rect 11227 8678 11279 8730
rect 11291 8678 11343 8730
rect 11355 8678 11407 8730
rect 31526 8678 31578 8730
rect 31590 8678 31642 8730
rect 31654 8678 31706 8730
rect 31718 8678 31770 8730
rect 51888 8678 51940 8730
rect 51952 8678 52004 8730
rect 52016 8678 52068 8730
rect 52080 8678 52132 8730
rect 2780 8576 2832 8628
rect 4068 8576 4120 8628
rect 5632 8576 5684 8628
rect 11520 8576 11572 8628
rect 3976 8440 4028 8492
rect 8392 8483 8444 8492
rect 1860 8415 1912 8424
rect 1860 8381 1869 8415
rect 1869 8381 1903 8415
rect 1903 8381 1912 8415
rect 1860 8372 1912 8381
rect 3148 8415 3200 8424
rect 3148 8381 3157 8415
rect 3157 8381 3191 8415
rect 3191 8381 3200 8415
rect 3148 8372 3200 8381
rect 5356 8415 5408 8424
rect 5356 8381 5365 8415
rect 5365 8381 5399 8415
rect 5399 8381 5408 8415
rect 5356 8372 5408 8381
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 14280 8576 14332 8628
rect 19432 8576 19484 8628
rect 13544 8551 13596 8560
rect 13544 8517 13553 8551
rect 13553 8517 13587 8551
rect 13587 8517 13596 8551
rect 13544 8508 13596 8517
rect 8668 8372 8720 8424
rect 10048 8372 10100 8424
rect 10876 8372 10928 8424
rect 11152 8415 11204 8424
rect 11152 8381 11161 8415
rect 11161 8381 11195 8415
rect 11195 8381 11204 8415
rect 11152 8372 11204 8381
rect 11612 8372 11664 8424
rect 13360 8372 13412 8424
rect 14648 8415 14700 8424
rect 14648 8381 14657 8415
rect 14657 8381 14691 8415
rect 14691 8381 14700 8415
rect 20720 8508 20772 8560
rect 21824 8576 21876 8628
rect 22008 8576 22060 8628
rect 32036 8576 32088 8628
rect 33048 8576 33100 8628
rect 34060 8576 34112 8628
rect 22192 8508 22244 8560
rect 22376 8508 22428 8560
rect 15568 8440 15620 8492
rect 20168 8440 20220 8492
rect 16028 8415 16080 8424
rect 14648 8372 14700 8381
rect 16028 8381 16037 8415
rect 16037 8381 16071 8415
rect 16071 8381 16080 8415
rect 18512 8415 18564 8424
rect 16028 8372 16080 8381
rect 18512 8381 18521 8415
rect 18521 8381 18555 8415
rect 18555 8381 18564 8415
rect 18512 8372 18564 8381
rect 18696 8415 18748 8424
rect 18696 8381 18705 8415
rect 18705 8381 18739 8415
rect 18739 8381 18748 8415
rect 18696 8372 18748 8381
rect 20076 8415 20128 8424
rect 17592 8304 17644 8356
rect 20076 8381 20085 8415
rect 20085 8381 20119 8415
rect 20119 8381 20128 8415
rect 20076 8372 20128 8381
rect 20536 8415 20588 8424
rect 20536 8381 20545 8415
rect 20545 8381 20579 8415
rect 20579 8381 20588 8415
rect 20536 8372 20588 8381
rect 20628 8415 20680 8424
rect 20628 8381 20637 8415
rect 20637 8381 20671 8415
rect 20671 8381 20680 8415
rect 20628 8372 20680 8381
rect 20812 8372 20864 8424
rect 22192 8372 22244 8424
rect 20904 8304 20956 8356
rect 21824 8304 21876 8356
rect 22468 8440 22520 8492
rect 23848 8551 23900 8560
rect 23848 8517 23857 8551
rect 23857 8517 23891 8551
rect 23891 8517 23900 8551
rect 23848 8508 23900 8517
rect 30840 8508 30892 8560
rect 36084 8576 36136 8628
rect 39304 8576 39356 8628
rect 39488 8619 39540 8628
rect 39488 8585 39497 8619
rect 39497 8585 39531 8619
rect 39531 8585 39540 8619
rect 39488 8576 39540 8585
rect 42064 8576 42116 8628
rect 44640 8576 44692 8628
rect 48136 8576 48188 8628
rect 50344 8576 50396 8628
rect 50436 8576 50488 8628
rect 52736 8619 52788 8628
rect 52736 8585 52745 8619
rect 52745 8585 52779 8619
rect 52779 8585 52788 8619
rect 52736 8576 52788 8585
rect 55036 8576 55088 8628
rect 58532 8576 58584 8628
rect 36544 8508 36596 8560
rect 37004 8508 37056 8560
rect 42156 8508 42208 8560
rect 42340 8508 42392 8560
rect 23388 8372 23440 8424
rect 24860 8372 24912 8424
rect 25412 8415 25464 8424
rect 25412 8381 25421 8415
rect 25421 8381 25455 8415
rect 25455 8381 25464 8415
rect 25412 8372 25464 8381
rect 26516 8440 26568 8492
rect 27804 8440 27856 8492
rect 30380 8440 30432 8492
rect 31852 8483 31904 8492
rect 31852 8449 31861 8483
rect 31861 8449 31895 8483
rect 31895 8449 31904 8483
rect 31852 8440 31904 8449
rect 33140 8440 33192 8492
rect 33876 8440 33928 8492
rect 34520 8440 34572 8492
rect 26884 8372 26936 8424
rect 27068 8372 27120 8424
rect 27436 8304 27488 8356
rect 27620 8347 27672 8356
rect 27620 8313 27629 8347
rect 27629 8313 27663 8347
rect 27663 8313 27672 8347
rect 27620 8304 27672 8313
rect 29552 8372 29604 8424
rect 29736 8415 29788 8424
rect 29736 8381 29745 8415
rect 29745 8381 29779 8415
rect 29779 8381 29788 8415
rect 29736 8372 29788 8381
rect 31024 8372 31076 8424
rect 32312 8372 32364 8424
rect 33232 8415 33284 8424
rect 33232 8381 33241 8415
rect 33241 8381 33275 8415
rect 33275 8381 33284 8415
rect 33232 8372 33284 8381
rect 33784 8415 33836 8424
rect 33784 8381 33793 8415
rect 33793 8381 33827 8415
rect 33827 8381 33836 8415
rect 33784 8372 33836 8381
rect 34888 8415 34940 8424
rect 34888 8381 34897 8415
rect 34897 8381 34931 8415
rect 34931 8381 34940 8415
rect 34888 8372 34940 8381
rect 35440 8415 35492 8424
rect 35440 8381 35449 8415
rect 35449 8381 35483 8415
rect 35483 8381 35492 8415
rect 35440 8372 35492 8381
rect 35716 8415 35768 8424
rect 35716 8381 35725 8415
rect 35725 8381 35759 8415
rect 35759 8381 35768 8415
rect 35716 8372 35768 8381
rect 36820 8415 36872 8424
rect 35624 8304 35676 8356
rect 36176 8304 36228 8356
rect 36820 8381 36829 8415
rect 36829 8381 36863 8415
rect 36863 8381 36872 8415
rect 36820 8372 36872 8381
rect 37280 8372 37332 8424
rect 38292 8372 38344 8424
rect 40040 8372 40092 8424
rect 41420 8372 41472 8424
rect 42156 8372 42208 8424
rect 42432 8372 42484 8424
rect 42800 8508 42852 8560
rect 46296 8508 46348 8560
rect 46940 8483 46992 8492
rect 46940 8449 46949 8483
rect 46949 8449 46983 8483
rect 46983 8449 46992 8483
rect 46940 8440 46992 8449
rect 42892 8372 42944 8424
rect 44180 8415 44232 8424
rect 44180 8381 44203 8415
rect 44203 8381 44232 8415
rect 44364 8415 44416 8424
rect 44180 8372 44232 8381
rect 44364 8381 44373 8415
rect 44373 8381 44407 8415
rect 44407 8381 44416 8415
rect 44364 8372 44416 8381
rect 44456 8372 44508 8424
rect 44824 8415 44876 8424
rect 44824 8381 44833 8415
rect 44833 8381 44867 8415
rect 44867 8381 44876 8415
rect 44824 8372 44876 8381
rect 45836 8415 45888 8424
rect 45836 8381 45845 8415
rect 45845 8381 45879 8415
rect 45879 8381 45888 8415
rect 45836 8372 45888 8381
rect 46296 8415 46348 8424
rect 46296 8381 46305 8415
rect 46305 8381 46339 8415
rect 46339 8381 46348 8415
rect 46296 8372 46348 8381
rect 46848 8415 46900 8424
rect 46848 8381 46857 8415
rect 46857 8381 46891 8415
rect 46891 8381 46900 8415
rect 46848 8372 46900 8381
rect 51356 8508 51408 8560
rect 48412 8440 48464 8492
rect 50252 8415 50304 8424
rect 50252 8381 50261 8415
rect 50261 8381 50295 8415
rect 50295 8381 50304 8415
rect 50252 8372 50304 8381
rect 50344 8415 50396 8424
rect 50344 8381 50353 8415
rect 50353 8381 50387 8415
rect 50387 8381 50396 8415
rect 50344 8372 50396 8381
rect 52184 8372 52236 8424
rect 53196 8415 53248 8424
rect 53196 8381 53219 8415
rect 53219 8381 53248 8415
rect 54944 8440 54996 8492
rect 55220 8508 55272 8560
rect 58808 8551 58860 8560
rect 58808 8517 58817 8551
rect 58817 8517 58851 8551
rect 58851 8517 58860 8551
rect 58808 8508 58860 8517
rect 59176 8440 59228 8492
rect 53196 8372 53248 8381
rect 53656 8415 53708 8424
rect 53656 8381 53665 8415
rect 53665 8381 53699 8415
rect 53699 8381 53708 8415
rect 53656 8372 53708 8381
rect 55864 8415 55916 8424
rect 46112 8304 46164 8356
rect 47952 8304 48004 8356
rect 55864 8381 55873 8415
rect 55873 8381 55907 8415
rect 55907 8381 55916 8415
rect 55864 8372 55916 8381
rect 56324 8372 56376 8424
rect 58532 8415 58584 8424
rect 58532 8381 58541 8415
rect 58541 8381 58575 8415
rect 58575 8381 58584 8415
rect 58532 8372 58584 8381
rect 59268 8415 59320 8424
rect 59268 8381 59277 8415
rect 59277 8381 59311 8415
rect 59311 8381 59320 8415
rect 59268 8372 59320 8381
rect 19984 8236 20036 8288
rect 20076 8236 20128 8288
rect 30656 8236 30708 8288
rect 32772 8236 32824 8288
rect 39764 8236 39816 8288
rect 40684 8279 40736 8288
rect 40684 8245 40693 8279
rect 40693 8245 40727 8279
rect 40727 8245 40736 8279
rect 40684 8236 40736 8245
rect 44824 8236 44876 8288
rect 45560 8236 45612 8288
rect 46020 8236 46072 8288
rect 46388 8236 46440 8288
rect 49608 8236 49660 8288
rect 50804 8236 50856 8288
rect 56876 8304 56928 8356
rect 56968 8304 57020 8356
rect 21344 8134 21396 8186
rect 21408 8134 21460 8186
rect 21472 8134 21524 8186
rect 21536 8134 21588 8186
rect 41707 8134 41759 8186
rect 41771 8134 41823 8186
rect 41835 8134 41887 8186
rect 41899 8134 41951 8186
rect 10784 8032 10836 8084
rect 2872 7896 2924 7948
rect 4068 7964 4120 8016
rect 4344 7964 4396 8016
rect 11152 7964 11204 8016
rect 3240 7896 3292 7948
rect 5080 7939 5132 7948
rect 5080 7905 5089 7939
rect 5089 7905 5123 7939
rect 5123 7905 5132 7939
rect 5080 7896 5132 7905
rect 3056 7871 3108 7880
rect 3056 7837 3065 7871
rect 3065 7837 3099 7871
rect 3099 7837 3108 7871
rect 5632 7896 5684 7948
rect 8300 7896 8352 7948
rect 10324 7939 10376 7948
rect 10324 7905 10333 7939
rect 10333 7905 10367 7939
rect 10367 7905 10376 7939
rect 10324 7896 10376 7905
rect 10692 7939 10744 7948
rect 10692 7905 10701 7939
rect 10701 7905 10735 7939
rect 10735 7905 10744 7939
rect 10692 7896 10744 7905
rect 15936 8032 15988 8084
rect 16488 8032 16540 8084
rect 17684 8032 17736 8084
rect 19708 8032 19760 8084
rect 22100 8032 22152 8084
rect 22192 8032 22244 8084
rect 12716 7964 12768 8016
rect 8760 7871 8812 7880
rect 3056 7828 3108 7837
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 12624 7896 12676 7948
rect 13544 7896 13596 7948
rect 13820 7828 13872 7880
rect 14648 7896 14700 7948
rect 16120 7896 16172 7948
rect 17592 7939 17644 7948
rect 17592 7905 17601 7939
rect 17601 7905 17635 7939
rect 17635 7905 17644 7939
rect 17592 7896 17644 7905
rect 17868 7964 17920 8016
rect 20444 7964 20496 8016
rect 20536 7964 20588 8016
rect 19524 7939 19576 7948
rect 15844 7828 15896 7880
rect 16580 7828 16632 7880
rect 18052 7828 18104 7880
rect 18696 7828 18748 7880
rect 19248 7828 19300 7880
rect 19524 7905 19533 7939
rect 19533 7905 19567 7939
rect 19567 7905 19576 7939
rect 19524 7896 19576 7905
rect 20628 7896 20680 7948
rect 20812 7896 20864 7948
rect 21088 7939 21140 7948
rect 21088 7905 21097 7939
rect 21097 7905 21131 7939
rect 21131 7905 21140 7939
rect 21088 7896 21140 7905
rect 22192 7896 22244 7948
rect 22560 7896 22612 7948
rect 23664 7896 23716 7948
rect 27344 7964 27396 8016
rect 27620 7964 27672 8016
rect 27160 7896 27212 7948
rect 27712 7896 27764 7948
rect 27804 7939 27856 7948
rect 27804 7905 27813 7939
rect 27813 7905 27847 7939
rect 27847 7905 27856 7939
rect 27804 7896 27856 7905
rect 27988 7939 28040 7948
rect 27988 7905 27997 7939
rect 27997 7905 28031 7939
rect 28031 7905 28040 7939
rect 29000 7939 29052 7948
rect 27988 7896 28040 7905
rect 29000 7905 29009 7939
rect 29009 7905 29043 7939
rect 29043 7905 29052 7939
rect 29000 7896 29052 7905
rect 20536 7828 20588 7880
rect 20720 7828 20772 7880
rect 22100 7828 22152 7880
rect 22284 7828 22336 7880
rect 22928 7828 22980 7880
rect 3148 7760 3200 7812
rect 6644 7760 6696 7812
rect 22468 7760 22520 7812
rect 27896 7828 27948 7880
rect 11796 7735 11848 7744
rect 11796 7701 11805 7735
rect 11805 7701 11839 7735
rect 11839 7701 11848 7735
rect 11796 7692 11848 7701
rect 14280 7735 14332 7744
rect 14280 7701 14289 7735
rect 14289 7701 14323 7735
rect 14323 7701 14332 7735
rect 14280 7692 14332 7701
rect 15384 7692 15436 7744
rect 15660 7692 15712 7744
rect 20352 7692 20404 7744
rect 25688 7692 25740 7744
rect 25780 7692 25832 7744
rect 31944 7964 31996 8016
rect 33232 7964 33284 8016
rect 33416 7964 33468 8016
rect 32036 7896 32088 7948
rect 32588 7939 32640 7948
rect 32588 7905 32597 7939
rect 32597 7905 32631 7939
rect 32631 7905 32640 7939
rect 32588 7896 32640 7905
rect 34520 7939 34572 7948
rect 34520 7905 34529 7939
rect 34529 7905 34563 7939
rect 34563 7905 34572 7939
rect 34520 7896 34572 7905
rect 34888 7939 34940 7948
rect 34888 7905 34897 7939
rect 34897 7905 34931 7939
rect 34931 7905 34940 7939
rect 34888 7896 34940 7905
rect 34980 7939 35032 7948
rect 34980 7905 34989 7939
rect 34989 7905 35023 7939
rect 35023 7905 35032 7939
rect 37372 7964 37424 8016
rect 39580 8007 39632 8016
rect 34980 7896 35032 7905
rect 36084 7939 36136 7948
rect 36084 7905 36093 7939
rect 36093 7905 36127 7939
rect 36127 7905 36136 7939
rect 36084 7896 36136 7905
rect 36268 7896 36320 7948
rect 37740 7939 37792 7948
rect 37740 7905 37749 7939
rect 37749 7905 37783 7939
rect 37783 7905 37792 7939
rect 37740 7896 37792 7905
rect 39304 7896 39356 7948
rect 31392 7828 31444 7880
rect 32404 7828 32456 7880
rect 33784 7828 33836 7880
rect 38844 7828 38896 7880
rect 39580 7973 39589 8007
rect 39589 7973 39623 8007
rect 39623 7973 39632 8007
rect 39580 7964 39632 7973
rect 39764 8032 39816 8084
rect 42340 7964 42392 8016
rect 40316 7896 40368 7948
rect 41236 7896 41288 7948
rect 41604 7896 41656 7948
rect 42248 7896 42300 7948
rect 43536 7896 43588 7948
rect 43996 7964 44048 8016
rect 44916 8032 44968 8084
rect 46112 8032 46164 8084
rect 46204 8032 46256 8084
rect 47768 8075 47820 8084
rect 47768 8041 47777 8075
rect 47777 8041 47811 8075
rect 47811 8041 47820 8075
rect 47768 8032 47820 8041
rect 55220 8075 55272 8084
rect 55220 8041 55229 8075
rect 55229 8041 55263 8075
rect 55263 8041 55272 8075
rect 55220 8032 55272 8041
rect 57244 8032 57296 8084
rect 44088 7939 44140 7948
rect 44088 7905 44097 7939
rect 44097 7905 44131 7939
rect 44131 7905 44140 7939
rect 44088 7896 44140 7905
rect 44456 7896 44508 7948
rect 51724 7964 51776 8016
rect 46112 7896 46164 7948
rect 47492 7896 47544 7948
rect 50436 7896 50488 7948
rect 51448 7939 51500 7948
rect 51448 7905 51457 7939
rect 51457 7905 51491 7939
rect 51491 7905 51500 7939
rect 51448 7896 51500 7905
rect 52460 7896 52512 7948
rect 55772 7964 55824 8016
rect 59268 7964 59320 8016
rect 55036 7939 55088 7948
rect 55036 7905 55045 7939
rect 55045 7905 55079 7939
rect 55079 7905 55088 7939
rect 55036 7896 55088 7905
rect 55312 7896 55364 7948
rect 56968 7939 57020 7948
rect 56968 7905 56977 7939
rect 56977 7905 57011 7939
rect 57011 7905 57020 7939
rect 56968 7896 57020 7905
rect 44732 7828 44784 7880
rect 45284 7828 45336 7880
rect 45560 7828 45612 7880
rect 45744 7828 45796 7880
rect 49792 7828 49844 7880
rect 50804 7871 50856 7880
rect 50804 7837 50813 7871
rect 50813 7837 50847 7871
rect 50847 7837 50856 7871
rect 50804 7828 50856 7837
rect 53104 7871 53156 7880
rect 53104 7837 53113 7871
rect 53113 7837 53147 7871
rect 53147 7837 53156 7871
rect 53104 7828 53156 7837
rect 55404 7828 55456 7880
rect 55680 7828 55732 7880
rect 60280 7939 60332 7948
rect 57244 7871 57296 7880
rect 57244 7837 57253 7871
rect 57253 7837 57287 7871
rect 57287 7837 57296 7871
rect 57244 7828 57296 7837
rect 57980 7828 58032 7880
rect 60280 7905 60289 7939
rect 60289 7905 60323 7939
rect 60323 7905 60332 7939
rect 60280 7896 60332 7905
rect 59452 7828 59504 7880
rect 32312 7692 32364 7744
rect 33600 7760 33652 7812
rect 42156 7803 42208 7812
rect 37096 7692 37148 7744
rect 38016 7692 38068 7744
rect 40408 7692 40460 7744
rect 42156 7769 42165 7803
rect 42165 7769 42199 7803
rect 42199 7769 42208 7803
rect 42156 7760 42208 7769
rect 43444 7735 43496 7744
rect 43444 7701 43453 7735
rect 43453 7701 43487 7735
rect 43487 7701 43496 7735
rect 43444 7692 43496 7701
rect 43536 7692 43588 7744
rect 51264 7760 51316 7812
rect 53748 7760 53800 7812
rect 54852 7803 54904 7812
rect 54852 7769 54861 7803
rect 54861 7769 54895 7803
rect 54895 7769 54904 7803
rect 54852 7760 54904 7769
rect 47216 7692 47268 7744
rect 58348 7735 58400 7744
rect 58348 7701 58357 7735
rect 58357 7701 58391 7735
rect 58391 7701 58400 7735
rect 58348 7692 58400 7701
rect 58808 7735 58860 7744
rect 58808 7701 58817 7735
rect 58817 7701 58851 7735
rect 58851 7701 58860 7735
rect 58808 7692 58860 7701
rect 60464 7735 60516 7744
rect 60464 7701 60473 7735
rect 60473 7701 60507 7735
rect 60507 7701 60516 7735
rect 60464 7692 60516 7701
rect 11163 7590 11215 7642
rect 11227 7590 11279 7642
rect 11291 7590 11343 7642
rect 11355 7590 11407 7642
rect 31526 7590 31578 7642
rect 31590 7590 31642 7642
rect 31654 7590 31706 7642
rect 31718 7590 31770 7642
rect 51888 7590 51940 7642
rect 51952 7590 52004 7642
rect 52016 7590 52068 7642
rect 52080 7590 52132 7642
rect 5632 7531 5684 7540
rect 5632 7497 5641 7531
rect 5641 7497 5675 7531
rect 5675 7497 5684 7531
rect 5632 7488 5684 7497
rect 13728 7488 13780 7540
rect 14924 7488 14976 7540
rect 9772 7420 9824 7472
rect 19524 7488 19576 7540
rect 19984 7488 20036 7540
rect 3976 7352 4028 7404
rect 8116 7352 8168 7404
rect 8668 7352 8720 7404
rect 8760 7352 8812 7404
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 4252 7216 4304 7268
rect 6644 7284 6696 7336
rect 9680 7284 9732 7336
rect 10968 7284 11020 7336
rect 12992 7352 13044 7404
rect 15016 7395 15068 7404
rect 9956 7259 10008 7268
rect 9956 7225 9965 7259
rect 9965 7225 9999 7259
rect 9999 7225 10008 7259
rect 13360 7284 13412 7336
rect 13452 7327 13504 7336
rect 13452 7293 13461 7327
rect 13461 7293 13495 7327
rect 13495 7293 13504 7327
rect 13452 7284 13504 7293
rect 14464 7327 14516 7336
rect 14464 7293 14473 7327
rect 14473 7293 14507 7327
rect 14507 7293 14516 7327
rect 14464 7284 14516 7293
rect 14648 7284 14700 7336
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 16488 7352 16540 7404
rect 17132 7395 17184 7404
rect 15936 7284 15988 7336
rect 16764 7284 16816 7336
rect 17132 7361 17141 7395
rect 17141 7361 17175 7395
rect 17175 7361 17184 7395
rect 17132 7352 17184 7361
rect 20076 7352 20128 7404
rect 18788 7327 18840 7336
rect 18788 7293 18797 7327
rect 18797 7293 18831 7327
rect 18831 7293 18840 7327
rect 18788 7284 18840 7293
rect 9956 7216 10008 7225
rect 11888 7216 11940 7268
rect 17960 7216 18012 7268
rect 4436 7191 4488 7200
rect 4436 7157 4445 7191
rect 4445 7157 4479 7191
rect 4479 7157 4488 7191
rect 4436 7148 4488 7157
rect 13452 7148 13504 7200
rect 15660 7148 15712 7200
rect 15752 7148 15804 7200
rect 16396 7148 16448 7200
rect 19708 7148 19760 7200
rect 20352 7420 20404 7472
rect 20628 7352 20680 7404
rect 21916 7352 21968 7404
rect 22284 7420 22336 7472
rect 25780 7463 25832 7472
rect 25780 7429 25789 7463
rect 25789 7429 25823 7463
rect 25823 7429 25832 7463
rect 25780 7420 25832 7429
rect 27988 7420 28040 7472
rect 31392 7420 31444 7472
rect 31944 7463 31996 7472
rect 31944 7429 31953 7463
rect 31953 7429 31987 7463
rect 31987 7429 31996 7463
rect 31944 7420 31996 7429
rect 32496 7488 32548 7540
rect 40316 7420 40368 7472
rect 44088 7488 44140 7540
rect 22008 7327 22060 7336
rect 20904 7216 20956 7268
rect 22008 7293 22017 7327
rect 22017 7293 22051 7327
rect 22051 7293 22060 7327
rect 22008 7284 22060 7293
rect 24216 7327 24268 7336
rect 24216 7293 24225 7327
rect 24225 7293 24259 7327
rect 24259 7293 24268 7327
rect 24216 7284 24268 7293
rect 22468 7216 22520 7268
rect 23296 7216 23348 7268
rect 25044 7216 25096 7268
rect 27160 7284 27212 7336
rect 27436 7284 27488 7336
rect 29000 7284 29052 7336
rect 29552 7284 29604 7336
rect 32864 7352 32916 7404
rect 33600 7395 33652 7404
rect 33600 7361 33609 7395
rect 33609 7361 33643 7395
rect 33643 7361 33652 7395
rect 33600 7352 33652 7361
rect 33784 7352 33836 7404
rect 36360 7352 36412 7404
rect 32588 7284 32640 7336
rect 33232 7327 33284 7336
rect 33232 7293 33241 7327
rect 33241 7293 33275 7327
rect 33275 7293 33284 7327
rect 33232 7284 33284 7293
rect 34336 7284 34388 7336
rect 35532 7327 35584 7336
rect 35532 7293 35541 7327
rect 35541 7293 35575 7327
rect 35575 7293 35584 7327
rect 35532 7284 35584 7293
rect 36084 7327 36136 7336
rect 36084 7293 36093 7327
rect 36093 7293 36127 7327
rect 36127 7293 36136 7327
rect 36084 7284 36136 7293
rect 36176 7284 36228 7336
rect 38108 7352 38160 7404
rect 38568 7352 38620 7404
rect 37004 7327 37056 7336
rect 37004 7293 37013 7327
rect 37013 7293 37047 7327
rect 37047 7293 37056 7327
rect 37004 7284 37056 7293
rect 37096 7284 37148 7336
rect 40684 7352 40736 7404
rect 42892 7352 42944 7404
rect 44272 7352 44324 7404
rect 44732 7395 44784 7404
rect 44732 7361 44741 7395
rect 44741 7361 44775 7395
rect 44775 7361 44784 7395
rect 44732 7352 44784 7361
rect 42156 7327 42208 7336
rect 42156 7293 42165 7327
rect 42165 7293 42199 7327
rect 42199 7293 42208 7327
rect 43076 7327 43128 7336
rect 42156 7284 42208 7293
rect 43076 7293 43085 7327
rect 43085 7293 43119 7327
rect 43119 7293 43128 7327
rect 43076 7284 43128 7293
rect 43996 7284 44048 7336
rect 46388 7352 46440 7404
rect 45192 7327 45244 7336
rect 45192 7293 45201 7327
rect 45201 7293 45235 7327
rect 45235 7293 45244 7327
rect 45192 7284 45244 7293
rect 46204 7284 46256 7336
rect 47492 7420 47544 7472
rect 47216 7352 47268 7404
rect 54760 7352 54812 7404
rect 56968 7352 57020 7404
rect 58072 7352 58124 7404
rect 58440 7352 58492 7404
rect 33048 7216 33100 7268
rect 35348 7216 35400 7268
rect 37280 7216 37332 7268
rect 38752 7216 38804 7268
rect 25596 7148 25648 7200
rect 29000 7148 29052 7200
rect 30472 7148 30524 7200
rect 30840 7191 30892 7200
rect 30840 7157 30849 7191
rect 30849 7157 30883 7191
rect 30883 7157 30892 7191
rect 30840 7148 30892 7157
rect 33784 7148 33836 7200
rect 35440 7148 35492 7200
rect 38568 7148 38620 7200
rect 41328 7216 41380 7268
rect 43352 7216 43404 7268
rect 46112 7259 46164 7268
rect 46112 7225 46121 7259
rect 46121 7225 46155 7259
rect 46155 7225 46164 7259
rect 46112 7216 46164 7225
rect 51540 7284 51592 7336
rect 51724 7284 51776 7336
rect 52552 7327 52604 7336
rect 52552 7293 52561 7327
rect 52561 7293 52595 7327
rect 52595 7293 52604 7327
rect 52552 7284 52604 7293
rect 55772 7327 55824 7336
rect 55772 7293 55781 7327
rect 55781 7293 55815 7327
rect 55815 7293 55824 7327
rect 55772 7284 55824 7293
rect 55864 7284 55916 7336
rect 50436 7216 50488 7268
rect 53932 7259 53984 7268
rect 53932 7225 53941 7259
rect 53941 7225 53975 7259
rect 53975 7225 53984 7259
rect 53932 7216 53984 7225
rect 54760 7216 54812 7268
rect 58624 7284 58676 7336
rect 42156 7148 42208 7200
rect 44732 7148 44784 7200
rect 47216 7148 47268 7200
rect 48228 7148 48280 7200
rect 53196 7148 53248 7200
rect 56968 7148 57020 7200
rect 59912 7191 59964 7200
rect 59912 7157 59921 7191
rect 59921 7157 59955 7191
rect 59955 7157 59964 7191
rect 59912 7148 59964 7157
rect 21344 7046 21396 7098
rect 21408 7046 21460 7098
rect 21472 7046 21524 7098
rect 21536 7046 21588 7098
rect 41707 7046 41759 7098
rect 41771 7046 41823 7098
rect 41835 7046 41887 7098
rect 41899 7046 41951 7098
rect 3056 6987 3108 6996
rect 3056 6953 3065 6987
rect 3065 6953 3099 6987
rect 3099 6953 3108 6987
rect 3056 6944 3108 6953
rect 3976 6808 4028 6860
rect 4160 6808 4212 6860
rect 5724 6851 5776 6860
rect 5724 6817 5733 6851
rect 5733 6817 5767 6851
rect 5767 6817 5776 6851
rect 5724 6808 5776 6817
rect 6460 6808 6512 6860
rect 6644 6851 6696 6860
rect 6644 6817 6653 6851
rect 6653 6817 6687 6851
rect 6687 6817 6696 6851
rect 6644 6808 6696 6817
rect 8760 6876 8812 6928
rect 8576 6851 8628 6860
rect 8576 6817 8585 6851
rect 8585 6817 8619 6851
rect 8619 6817 8628 6851
rect 10048 6876 10100 6928
rect 16120 6876 16172 6928
rect 18052 6876 18104 6928
rect 18788 6876 18840 6928
rect 8576 6808 8628 6817
rect 9956 6808 10008 6860
rect 10600 6851 10652 6860
rect 10600 6817 10609 6851
rect 10609 6817 10643 6851
rect 10643 6817 10652 6851
rect 10600 6808 10652 6817
rect 11888 6851 11940 6860
rect 11888 6817 11897 6851
rect 11897 6817 11931 6851
rect 11931 6817 11940 6851
rect 11888 6808 11940 6817
rect 12164 6808 12216 6860
rect 13820 6851 13872 6860
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 4344 6740 4396 6749
rect 7748 6740 7800 6792
rect 10324 6740 10376 6792
rect 11980 6783 12032 6792
rect 11980 6749 11989 6783
rect 11989 6749 12023 6783
rect 12023 6749 12032 6783
rect 11980 6740 12032 6749
rect 10140 6715 10192 6724
rect 10140 6681 10149 6715
rect 10149 6681 10183 6715
rect 10183 6681 10192 6715
rect 10140 6672 10192 6681
rect 13820 6817 13829 6851
rect 13829 6817 13863 6851
rect 13863 6817 13872 6851
rect 13820 6808 13872 6817
rect 14096 6808 14148 6860
rect 15108 6808 15160 6860
rect 20260 6876 20312 6928
rect 13084 6740 13136 6792
rect 19708 6851 19760 6860
rect 19708 6817 19717 6851
rect 19717 6817 19751 6851
rect 19751 6817 19760 6851
rect 19708 6808 19760 6817
rect 20904 6851 20956 6860
rect 20904 6817 20913 6851
rect 20913 6817 20947 6851
rect 20947 6817 20956 6851
rect 20904 6808 20956 6817
rect 20996 6808 21048 6860
rect 23388 6851 23440 6860
rect 15752 6740 15804 6792
rect 16304 6783 16356 6792
rect 16304 6749 16313 6783
rect 16313 6749 16347 6783
rect 16347 6749 16356 6783
rect 16304 6740 16356 6749
rect 19248 6783 19300 6792
rect 19248 6749 19257 6783
rect 19257 6749 19291 6783
rect 19291 6749 19300 6783
rect 19248 6740 19300 6749
rect 19524 6740 19576 6792
rect 22376 6740 22428 6792
rect 23388 6817 23397 6851
rect 23397 6817 23431 6851
rect 23431 6817 23440 6851
rect 23388 6808 23440 6817
rect 23572 6808 23624 6860
rect 25044 6851 25096 6860
rect 25044 6817 25053 6851
rect 25053 6817 25087 6851
rect 25087 6817 25096 6851
rect 25044 6808 25096 6817
rect 25688 6876 25740 6928
rect 27160 6919 27212 6928
rect 27160 6885 27169 6919
rect 27169 6885 27203 6919
rect 27203 6885 27212 6919
rect 27160 6876 27212 6885
rect 37188 6944 37240 6996
rect 37740 6944 37792 6996
rect 45560 6944 45612 6996
rect 23848 6740 23900 6792
rect 26884 6808 26936 6860
rect 26976 6851 27028 6860
rect 26976 6817 26985 6851
rect 26985 6817 27019 6851
rect 27019 6817 27028 6851
rect 26976 6808 27028 6817
rect 27804 6808 27856 6860
rect 27988 6851 28040 6860
rect 27988 6817 27997 6851
rect 27997 6817 28031 6851
rect 28031 6817 28040 6851
rect 27988 6808 28040 6817
rect 28080 6851 28132 6860
rect 28080 6817 28089 6851
rect 28089 6817 28123 6851
rect 28123 6817 28132 6851
rect 28080 6808 28132 6817
rect 28264 6808 28316 6860
rect 25964 6740 26016 6792
rect 14464 6672 14516 6724
rect 17960 6672 18012 6724
rect 25228 6672 25280 6724
rect 27528 6672 27580 6724
rect 28540 6808 28592 6860
rect 28724 6740 28776 6792
rect 30564 6808 30616 6860
rect 30656 6808 30708 6860
rect 32312 6808 32364 6860
rect 32680 6851 32732 6860
rect 32680 6817 32689 6851
rect 32689 6817 32723 6851
rect 32723 6817 32732 6851
rect 32680 6808 32732 6817
rect 33416 6808 33468 6860
rect 41236 6876 41288 6928
rect 33784 6851 33836 6860
rect 33784 6817 33793 6851
rect 33793 6817 33827 6851
rect 33827 6817 33836 6851
rect 33784 6808 33836 6817
rect 34888 6808 34940 6860
rect 35532 6808 35584 6860
rect 35992 6851 36044 6860
rect 35992 6817 36001 6851
rect 36001 6817 36035 6851
rect 36035 6817 36044 6851
rect 35992 6808 36044 6817
rect 36176 6851 36228 6860
rect 36176 6817 36185 6851
rect 36185 6817 36219 6851
rect 36219 6817 36228 6851
rect 36176 6808 36228 6817
rect 36360 6851 36412 6860
rect 36360 6817 36369 6851
rect 36369 6817 36403 6851
rect 36403 6817 36412 6851
rect 36360 6808 36412 6817
rect 36452 6808 36504 6860
rect 37004 6808 37056 6860
rect 37556 6808 37608 6860
rect 37740 6851 37792 6860
rect 37740 6817 37749 6851
rect 37749 6817 37783 6851
rect 37783 6817 37792 6851
rect 37740 6808 37792 6817
rect 38200 6808 38252 6860
rect 38752 6851 38804 6860
rect 38752 6817 38761 6851
rect 38761 6817 38795 6851
rect 38795 6817 38804 6851
rect 38752 6808 38804 6817
rect 38936 6851 38988 6860
rect 38936 6817 38945 6851
rect 38945 6817 38979 6851
rect 38979 6817 38988 6851
rect 38936 6808 38988 6817
rect 40408 6851 40460 6860
rect 40408 6817 40417 6851
rect 40417 6817 40451 6851
rect 40451 6817 40460 6851
rect 40868 6851 40920 6860
rect 40408 6808 40460 6817
rect 40868 6817 40877 6851
rect 40877 6817 40911 6851
rect 40911 6817 40920 6851
rect 40868 6808 40920 6817
rect 32496 6672 32548 6724
rect 32864 6715 32916 6724
rect 32864 6681 32873 6715
rect 32873 6681 32907 6715
rect 32907 6681 32916 6715
rect 32864 6672 32916 6681
rect 5540 6604 5592 6656
rect 10232 6604 10284 6656
rect 13084 6604 13136 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 19340 6604 19392 6656
rect 20260 6604 20312 6656
rect 26608 6604 26660 6656
rect 29460 6604 29512 6656
rect 30012 6647 30064 6656
rect 30012 6613 30021 6647
rect 30021 6613 30055 6647
rect 30055 6613 30064 6647
rect 30012 6604 30064 6613
rect 30104 6604 30156 6656
rect 41604 6740 41656 6792
rect 41972 6851 42024 6860
rect 41972 6817 41981 6851
rect 41981 6817 42015 6851
rect 42015 6817 42024 6851
rect 41972 6808 42024 6817
rect 42708 6808 42760 6860
rect 43904 6851 43956 6860
rect 43904 6817 43913 6851
rect 43913 6817 43947 6851
rect 43947 6817 43956 6851
rect 43904 6808 43956 6817
rect 44272 6808 44324 6860
rect 33324 6672 33376 6724
rect 41052 6672 41104 6724
rect 43444 6740 43496 6792
rect 44364 6783 44416 6792
rect 44364 6749 44373 6783
rect 44373 6749 44407 6783
rect 44407 6749 44416 6783
rect 44364 6740 44416 6749
rect 44916 6740 44968 6792
rect 45652 6808 45704 6860
rect 46756 6851 46808 6860
rect 46756 6817 46765 6851
rect 46765 6817 46799 6851
rect 46799 6817 46808 6851
rect 46756 6808 46808 6817
rect 47032 6851 47084 6860
rect 47032 6817 47041 6851
rect 47041 6817 47075 6851
rect 47075 6817 47084 6851
rect 47032 6808 47084 6817
rect 51356 6876 51408 6928
rect 52552 6876 52604 6928
rect 46112 6740 46164 6792
rect 46572 6740 46624 6792
rect 47308 6783 47360 6792
rect 47308 6749 47317 6783
rect 47317 6749 47351 6783
rect 47351 6749 47360 6783
rect 47308 6740 47360 6749
rect 48688 6740 48740 6792
rect 51264 6808 51316 6860
rect 53196 6876 53248 6928
rect 53656 6876 53708 6928
rect 49332 6740 49384 6792
rect 49516 6783 49568 6792
rect 49516 6749 49525 6783
rect 49525 6749 49559 6783
rect 49559 6749 49568 6783
rect 49516 6740 49568 6749
rect 46848 6715 46900 6724
rect 46848 6681 46857 6715
rect 46857 6681 46891 6715
rect 46891 6681 46900 6715
rect 46848 6672 46900 6681
rect 52368 6740 52420 6792
rect 53288 6740 53340 6792
rect 33232 6604 33284 6656
rect 39488 6604 39540 6656
rect 42616 6604 42668 6656
rect 52184 6672 52236 6724
rect 53840 6808 53892 6860
rect 54760 6851 54812 6860
rect 54760 6817 54769 6851
rect 54769 6817 54803 6851
rect 54803 6817 54812 6851
rect 54760 6808 54812 6817
rect 47032 6604 47084 6656
rect 47952 6604 48004 6656
rect 48044 6604 48096 6656
rect 51264 6604 51316 6656
rect 52920 6604 52972 6656
rect 53012 6604 53064 6656
rect 53748 6740 53800 6792
rect 56140 6808 56192 6860
rect 56692 6851 56744 6860
rect 56692 6817 56701 6851
rect 56701 6817 56735 6851
rect 56735 6817 56744 6851
rect 56692 6808 56744 6817
rect 58624 6876 58676 6928
rect 59360 6876 59412 6928
rect 56968 6851 57020 6860
rect 56968 6817 56977 6851
rect 56977 6817 57011 6851
rect 57011 6817 57020 6851
rect 56968 6808 57020 6817
rect 57980 6808 58032 6860
rect 58716 6851 58768 6860
rect 58716 6817 58725 6851
rect 58725 6817 58759 6851
rect 58759 6817 58768 6851
rect 58716 6808 58768 6817
rect 58808 6851 58860 6860
rect 58808 6817 58817 6851
rect 58817 6817 58851 6851
rect 58851 6817 58860 6851
rect 58808 6808 58860 6817
rect 56232 6783 56284 6792
rect 56232 6749 56241 6783
rect 56241 6749 56275 6783
rect 56275 6749 56284 6783
rect 59912 6808 59964 6860
rect 60280 6851 60332 6860
rect 60280 6817 60289 6851
rect 60289 6817 60323 6851
rect 60323 6817 60332 6851
rect 60280 6808 60332 6817
rect 56232 6740 56284 6749
rect 59544 6740 59596 6792
rect 60188 6783 60240 6792
rect 60188 6749 60197 6783
rect 60197 6749 60231 6783
rect 60231 6749 60240 6783
rect 60188 6740 60240 6749
rect 59268 6672 59320 6724
rect 54024 6604 54076 6656
rect 60280 6604 60332 6656
rect 11163 6502 11215 6554
rect 11227 6502 11279 6554
rect 11291 6502 11343 6554
rect 11355 6502 11407 6554
rect 31526 6502 31578 6554
rect 31590 6502 31642 6554
rect 31654 6502 31706 6554
rect 31718 6502 31770 6554
rect 51888 6502 51940 6554
rect 51952 6502 52004 6554
rect 52016 6502 52068 6554
rect 52080 6502 52132 6554
rect 9680 6443 9732 6452
rect 9680 6409 9689 6443
rect 9689 6409 9723 6443
rect 9723 6409 9732 6443
rect 9680 6400 9732 6409
rect 23572 6400 23624 6452
rect 3148 6264 3200 6316
rect 2688 6239 2740 6248
rect 2688 6205 2697 6239
rect 2697 6205 2731 6239
rect 2731 6205 2740 6239
rect 2688 6196 2740 6205
rect 5632 6264 5684 6316
rect 4436 6196 4488 6248
rect 4804 6196 4856 6248
rect 5356 6196 5408 6248
rect 17132 6332 17184 6384
rect 6368 6264 6420 6316
rect 10140 6307 10192 6316
rect 6920 6196 6972 6248
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 11980 6264 12032 6316
rect 12532 6264 12584 6316
rect 16212 6264 16264 6316
rect 16304 6264 16356 6316
rect 10232 6239 10284 6248
rect 10232 6205 10241 6239
rect 10241 6205 10275 6239
rect 10275 6205 10284 6239
rect 10232 6196 10284 6205
rect 10600 6239 10652 6248
rect 10600 6205 10609 6239
rect 10609 6205 10643 6239
rect 10643 6205 10652 6239
rect 10600 6196 10652 6205
rect 2780 6103 2832 6112
rect 2780 6069 2789 6103
rect 2789 6069 2823 6103
rect 2823 6069 2832 6103
rect 12532 6128 12584 6180
rect 15016 6171 15068 6180
rect 15016 6137 15025 6171
rect 15025 6137 15059 6171
rect 15059 6137 15068 6171
rect 15016 6128 15068 6137
rect 15476 6196 15528 6248
rect 16580 6196 16632 6248
rect 19892 6332 19944 6384
rect 20076 6332 20128 6384
rect 20168 6332 20220 6384
rect 19524 6307 19576 6316
rect 19524 6273 19533 6307
rect 19533 6273 19567 6307
rect 19567 6273 19576 6307
rect 19524 6264 19576 6273
rect 20720 6264 20772 6316
rect 27804 6332 27856 6384
rect 28264 6400 28316 6452
rect 33232 6400 33284 6452
rect 28356 6332 28408 6384
rect 36176 6400 36228 6452
rect 36912 6400 36964 6452
rect 38844 6400 38896 6452
rect 40684 6400 40736 6452
rect 41972 6400 42024 6452
rect 42340 6400 42392 6452
rect 48320 6400 48372 6452
rect 35992 6332 36044 6384
rect 36452 6332 36504 6384
rect 36820 6332 36872 6384
rect 38936 6332 38988 6384
rect 39672 6332 39724 6384
rect 49332 6332 49384 6384
rect 25228 6307 25280 6316
rect 20260 6239 20312 6248
rect 20260 6205 20269 6239
rect 20269 6205 20303 6239
rect 20303 6205 20312 6239
rect 20260 6196 20312 6205
rect 20352 6239 20404 6248
rect 20352 6205 20361 6239
rect 20361 6205 20395 6239
rect 20395 6205 20404 6239
rect 20352 6196 20404 6205
rect 20812 6196 20864 6248
rect 21548 6239 21600 6248
rect 21548 6205 21557 6239
rect 21557 6205 21591 6239
rect 21591 6205 21600 6239
rect 21548 6196 21600 6205
rect 21916 6196 21968 6248
rect 24952 6239 25004 6248
rect 22744 6128 22796 6180
rect 2780 6060 2832 6069
rect 7012 6060 7064 6112
rect 7104 6103 7156 6112
rect 7104 6069 7113 6103
rect 7113 6069 7147 6103
rect 7147 6069 7156 6103
rect 7104 6060 7156 6069
rect 7288 6060 7340 6112
rect 12072 6060 12124 6112
rect 12624 6103 12676 6112
rect 12624 6069 12633 6103
rect 12633 6069 12667 6103
rect 12667 6069 12676 6103
rect 12624 6060 12676 6069
rect 12716 6103 12768 6112
rect 12716 6069 12725 6103
rect 12725 6069 12759 6103
rect 12759 6069 12768 6103
rect 12716 6060 12768 6069
rect 16672 6060 16724 6112
rect 18696 6060 18748 6112
rect 21732 6103 21784 6112
rect 21732 6069 21741 6103
rect 21741 6069 21775 6103
rect 21775 6069 21784 6103
rect 21732 6060 21784 6069
rect 24032 6103 24084 6112
rect 24032 6069 24041 6103
rect 24041 6069 24075 6103
rect 24075 6069 24084 6103
rect 24032 6060 24084 6069
rect 24952 6205 24961 6239
rect 24961 6205 24995 6239
rect 24995 6205 25004 6239
rect 24952 6196 25004 6205
rect 25228 6273 25237 6307
rect 25237 6273 25271 6307
rect 25271 6273 25280 6307
rect 25228 6264 25280 6273
rect 33324 6264 33376 6316
rect 28908 6196 28960 6248
rect 29368 6196 29420 6248
rect 29460 6196 29512 6248
rect 31208 6196 31260 6248
rect 31300 6239 31352 6248
rect 31300 6205 31309 6239
rect 31309 6205 31343 6239
rect 31343 6205 31352 6239
rect 31300 6196 31352 6205
rect 30472 6128 30524 6180
rect 30932 6128 30984 6180
rect 31760 6196 31812 6248
rect 39396 6264 39448 6316
rect 41696 6264 41748 6316
rect 44916 6264 44968 6316
rect 34060 6196 34112 6248
rect 34244 6196 34296 6248
rect 36452 6239 36504 6248
rect 25964 6060 26016 6112
rect 29276 6060 29328 6112
rect 29460 6103 29512 6112
rect 29460 6069 29469 6103
rect 29469 6069 29503 6103
rect 29503 6069 29512 6103
rect 29460 6060 29512 6069
rect 30012 6060 30064 6112
rect 35900 6128 35952 6180
rect 35072 6103 35124 6112
rect 35072 6069 35081 6103
rect 35081 6069 35115 6103
rect 35115 6069 35124 6103
rect 35072 6060 35124 6069
rect 36452 6205 36461 6239
rect 36461 6205 36495 6239
rect 36495 6205 36504 6239
rect 36452 6196 36504 6205
rect 36912 6239 36964 6248
rect 36912 6205 36921 6239
rect 36921 6205 36955 6239
rect 36955 6205 36964 6239
rect 36912 6196 36964 6205
rect 37096 6196 37148 6248
rect 37648 6196 37700 6248
rect 39120 6239 39172 6248
rect 39120 6205 39129 6239
rect 39129 6205 39163 6239
rect 39163 6205 39172 6239
rect 39120 6196 39172 6205
rect 36360 6171 36412 6180
rect 36360 6137 36369 6171
rect 36369 6137 36403 6171
rect 36403 6137 36412 6171
rect 36360 6128 36412 6137
rect 39488 6128 39540 6180
rect 40408 6128 40460 6180
rect 40684 6239 40736 6248
rect 40684 6205 40693 6239
rect 40693 6205 40727 6239
rect 40727 6205 40736 6239
rect 40684 6196 40736 6205
rect 41420 6196 41472 6248
rect 42248 6196 42300 6248
rect 42616 6239 42668 6248
rect 42616 6205 42625 6239
rect 42625 6205 42659 6239
rect 42659 6205 42668 6239
rect 42616 6196 42668 6205
rect 42892 6239 42944 6248
rect 42892 6205 42901 6239
rect 42901 6205 42935 6239
rect 42935 6205 42944 6239
rect 42892 6196 42944 6205
rect 44640 6239 44692 6248
rect 44640 6205 44649 6239
rect 44649 6205 44683 6239
rect 44683 6205 44692 6239
rect 44640 6196 44692 6205
rect 53012 6400 53064 6452
rect 53564 6400 53616 6452
rect 53748 6400 53800 6452
rect 58164 6400 58216 6452
rect 49792 6332 49844 6384
rect 51632 6332 51684 6384
rect 52184 6332 52236 6384
rect 50528 6264 50580 6316
rect 51172 6264 51224 6316
rect 56692 6332 56744 6384
rect 53564 6264 53616 6316
rect 53932 6264 53984 6316
rect 54668 6264 54720 6316
rect 42340 6128 42392 6180
rect 42432 6128 42484 6180
rect 46296 6128 46348 6180
rect 48688 6239 48740 6248
rect 48688 6205 48697 6239
rect 48697 6205 48731 6239
rect 48731 6205 48740 6239
rect 48688 6196 48740 6205
rect 48872 6196 48924 6248
rect 49516 6196 49568 6248
rect 50620 6196 50672 6248
rect 51448 6196 51500 6248
rect 52828 6196 52880 6248
rect 53288 6196 53340 6248
rect 54484 6196 54536 6248
rect 54576 6239 54628 6248
rect 54576 6205 54585 6239
rect 54585 6205 54619 6239
rect 54619 6205 54628 6239
rect 55128 6239 55180 6248
rect 54576 6196 54628 6205
rect 55128 6205 55137 6239
rect 55137 6205 55171 6239
rect 55171 6205 55180 6239
rect 55128 6196 55180 6205
rect 55404 6239 55456 6248
rect 55404 6205 55413 6239
rect 55413 6205 55447 6239
rect 55447 6205 55456 6239
rect 55404 6196 55456 6205
rect 36452 6060 36504 6112
rect 42800 6060 42852 6112
rect 45560 6060 45612 6112
rect 49608 6128 49660 6180
rect 49792 6128 49844 6180
rect 53012 6171 53064 6180
rect 53012 6137 53021 6171
rect 53021 6137 53055 6171
rect 53055 6137 53064 6171
rect 53012 6128 53064 6137
rect 53748 6128 53800 6180
rect 58716 6239 58768 6248
rect 46756 6060 46808 6112
rect 50712 6060 50764 6112
rect 52184 6060 52236 6112
rect 56232 6060 56284 6112
rect 58716 6205 58725 6239
rect 58725 6205 58759 6239
rect 58759 6205 58768 6239
rect 58716 6196 58768 6205
rect 58808 6239 58860 6248
rect 58808 6205 58817 6239
rect 58817 6205 58851 6239
rect 58851 6205 58860 6239
rect 59268 6264 59320 6316
rect 58808 6196 58860 6205
rect 59176 6239 59228 6248
rect 59176 6205 59185 6239
rect 59185 6205 59219 6239
rect 59219 6205 59228 6239
rect 59544 6264 59596 6316
rect 59176 6196 59228 6205
rect 58072 6171 58124 6180
rect 58072 6137 58081 6171
rect 58081 6137 58115 6171
rect 58115 6137 58124 6171
rect 58072 6128 58124 6137
rect 57796 6060 57848 6112
rect 21344 5958 21396 6010
rect 21408 5958 21460 6010
rect 21472 5958 21524 6010
rect 21536 5958 21588 6010
rect 41707 5958 41759 6010
rect 41771 5958 41823 6010
rect 41835 5958 41887 6010
rect 41899 5958 41951 6010
rect 8208 5856 8260 5908
rect 8944 5856 8996 5908
rect 12716 5856 12768 5908
rect 13820 5856 13872 5908
rect 23204 5856 23256 5908
rect 27160 5856 27212 5908
rect 27252 5856 27304 5908
rect 30932 5856 30984 5908
rect 31300 5856 31352 5908
rect 35072 5856 35124 5908
rect 37924 5856 37976 5908
rect 39028 5856 39080 5908
rect 4344 5788 4396 5840
rect 4252 5720 4304 5772
rect 5540 5788 5592 5840
rect 4804 5763 4856 5772
rect 4804 5729 4813 5763
rect 4813 5729 4847 5763
rect 4847 5729 4856 5763
rect 4804 5720 4856 5729
rect 5724 5720 5776 5772
rect 6736 5788 6788 5840
rect 15016 5788 15068 5840
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 2872 5516 2924 5525
rect 7288 5720 7340 5772
rect 7932 5763 7984 5772
rect 7932 5729 7941 5763
rect 7941 5729 7975 5763
rect 7975 5729 7984 5763
rect 7932 5720 7984 5729
rect 8024 5720 8076 5772
rect 11796 5720 11848 5772
rect 12348 5720 12400 5772
rect 12440 5720 12492 5772
rect 15200 5720 15252 5772
rect 15660 5763 15712 5772
rect 15660 5729 15669 5763
rect 15669 5729 15703 5763
rect 15703 5729 15712 5763
rect 15660 5720 15712 5729
rect 15752 5720 15804 5772
rect 16396 5720 16448 5772
rect 21180 5788 21232 5840
rect 23480 5788 23532 5840
rect 25596 5788 25648 5840
rect 19340 5763 19392 5772
rect 19340 5729 19349 5763
rect 19349 5729 19383 5763
rect 19383 5729 19392 5763
rect 19340 5720 19392 5729
rect 21088 5720 21140 5772
rect 24860 5763 24912 5772
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 12532 5652 12584 5704
rect 12624 5652 12676 5704
rect 15384 5652 15436 5704
rect 16304 5652 16356 5704
rect 20076 5652 20128 5704
rect 24860 5729 24869 5763
rect 24869 5729 24903 5763
rect 24903 5729 24912 5763
rect 24860 5720 24912 5729
rect 25228 5763 25280 5772
rect 25228 5729 25237 5763
rect 25237 5729 25271 5763
rect 25271 5729 25280 5763
rect 25228 5720 25280 5729
rect 25320 5720 25372 5772
rect 26976 5763 27028 5772
rect 26976 5729 26985 5763
rect 26985 5729 27019 5763
rect 27019 5729 27028 5763
rect 26976 5720 27028 5729
rect 27252 5720 27304 5772
rect 27988 5788 28040 5840
rect 28356 5788 28408 5840
rect 27528 5720 27580 5772
rect 27712 5720 27764 5772
rect 30196 5788 30248 5840
rect 32404 5788 32456 5840
rect 34612 5788 34664 5840
rect 39120 5788 39172 5840
rect 39488 5788 39540 5840
rect 42800 5856 42852 5908
rect 42892 5856 42944 5908
rect 30104 5720 30156 5772
rect 30932 5720 30984 5772
rect 31116 5720 31168 5772
rect 32312 5763 32364 5772
rect 32312 5729 32321 5763
rect 32321 5729 32355 5763
rect 32355 5729 32364 5763
rect 32312 5720 32364 5729
rect 32588 5720 32640 5772
rect 37188 5720 37240 5772
rect 38752 5720 38804 5772
rect 39396 5763 39448 5772
rect 39396 5729 39405 5763
rect 39405 5729 39439 5763
rect 39439 5729 39448 5763
rect 39396 5720 39448 5729
rect 40868 5763 40920 5772
rect 40868 5729 40877 5763
rect 40877 5729 40911 5763
rect 40911 5729 40920 5763
rect 44640 5788 44692 5840
rect 40868 5720 40920 5729
rect 42340 5720 42392 5772
rect 44088 5720 44140 5772
rect 44456 5763 44508 5772
rect 44456 5729 44465 5763
rect 44465 5729 44499 5763
rect 44499 5729 44508 5763
rect 44456 5720 44508 5729
rect 47216 5856 47268 5908
rect 48872 5856 48924 5908
rect 49424 5899 49476 5908
rect 49424 5865 49433 5899
rect 49433 5865 49467 5899
rect 49467 5865 49476 5899
rect 49424 5856 49476 5865
rect 49884 5788 49936 5840
rect 50252 5856 50304 5908
rect 50528 5856 50580 5908
rect 52460 5856 52512 5908
rect 50620 5788 50672 5840
rect 51540 5831 51592 5840
rect 51540 5797 51549 5831
rect 51549 5797 51583 5831
rect 51583 5797 51592 5831
rect 51540 5788 51592 5797
rect 52828 5856 52880 5908
rect 45652 5763 45704 5772
rect 45652 5729 45661 5763
rect 45661 5729 45695 5763
rect 45695 5729 45704 5763
rect 45652 5720 45704 5729
rect 6920 5627 6972 5636
rect 6920 5593 6929 5627
rect 6929 5593 6963 5627
rect 6963 5593 6972 5627
rect 6920 5584 6972 5593
rect 10968 5584 11020 5636
rect 15292 5584 15344 5636
rect 22376 5584 22428 5636
rect 29276 5652 29328 5704
rect 30196 5695 30248 5704
rect 30196 5661 30205 5695
rect 30205 5661 30239 5695
rect 30239 5661 30248 5695
rect 30196 5652 30248 5661
rect 30472 5652 30524 5704
rect 32680 5695 32732 5704
rect 32680 5661 32689 5695
rect 32689 5661 32723 5695
rect 32723 5661 32732 5695
rect 32680 5652 32732 5661
rect 33232 5652 33284 5704
rect 34060 5652 34112 5704
rect 34336 5695 34388 5704
rect 34336 5661 34345 5695
rect 34345 5661 34379 5695
rect 34379 5661 34388 5695
rect 34336 5652 34388 5661
rect 26424 5584 26476 5636
rect 27712 5584 27764 5636
rect 12440 5559 12492 5568
rect 12440 5525 12449 5559
rect 12449 5525 12483 5559
rect 12483 5525 12492 5559
rect 13728 5559 13780 5568
rect 12440 5516 12492 5525
rect 13728 5525 13737 5559
rect 13737 5525 13771 5559
rect 13771 5525 13780 5559
rect 13728 5516 13780 5525
rect 15476 5516 15528 5568
rect 17500 5516 17552 5568
rect 17960 5516 18012 5568
rect 19340 5516 19392 5568
rect 23112 5559 23164 5568
rect 23112 5525 23121 5559
rect 23121 5525 23155 5559
rect 23155 5525 23164 5559
rect 23112 5516 23164 5525
rect 23572 5559 23624 5568
rect 23572 5525 23581 5559
rect 23581 5525 23615 5559
rect 23615 5525 23624 5559
rect 23572 5516 23624 5525
rect 23848 5516 23900 5568
rect 28816 5516 28868 5568
rect 29092 5559 29144 5568
rect 29092 5525 29101 5559
rect 29101 5525 29135 5559
rect 29135 5525 29144 5559
rect 29092 5516 29144 5525
rect 31852 5584 31904 5636
rect 45192 5652 45244 5704
rect 45468 5695 45520 5704
rect 45468 5661 45477 5695
rect 45477 5661 45511 5695
rect 45511 5661 45520 5695
rect 45468 5652 45520 5661
rect 34520 5584 34572 5636
rect 36176 5584 36228 5636
rect 36360 5584 36412 5636
rect 46388 5652 46440 5704
rect 48044 5695 48096 5704
rect 45652 5584 45704 5636
rect 47216 5584 47268 5636
rect 48044 5661 48053 5695
rect 48053 5661 48087 5695
rect 48087 5661 48096 5695
rect 48044 5652 48096 5661
rect 48136 5652 48188 5704
rect 49240 5695 49292 5704
rect 49240 5661 49249 5695
rect 49249 5661 49283 5695
rect 49283 5661 49292 5695
rect 49240 5652 49292 5661
rect 50436 5720 50488 5772
rect 51264 5720 51316 5772
rect 56508 5856 56560 5908
rect 57520 5856 57572 5908
rect 53472 5788 53524 5840
rect 55404 5788 55456 5840
rect 49792 5652 49844 5704
rect 47676 5584 47728 5636
rect 52092 5720 52144 5772
rect 53380 5720 53432 5772
rect 57796 5763 57848 5772
rect 36268 5516 36320 5568
rect 37280 5516 37332 5568
rect 40592 5559 40644 5568
rect 40592 5525 40601 5559
rect 40601 5525 40635 5559
rect 40635 5525 40644 5559
rect 40592 5516 40644 5525
rect 42064 5516 42116 5568
rect 42432 5516 42484 5568
rect 52092 5584 52144 5636
rect 52368 5584 52420 5636
rect 54760 5652 54812 5704
rect 56232 5652 56284 5704
rect 57796 5729 57805 5763
rect 57805 5729 57839 5763
rect 57839 5729 57848 5763
rect 57796 5720 57848 5729
rect 59176 5788 59228 5840
rect 57520 5652 57572 5704
rect 53840 5584 53892 5636
rect 54392 5584 54444 5636
rect 52276 5516 52328 5568
rect 56324 5516 56376 5568
rect 57704 5584 57756 5636
rect 58348 5516 58400 5568
rect 58624 5516 58676 5568
rect 58808 5516 58860 5568
rect 11163 5414 11215 5466
rect 11227 5414 11279 5466
rect 11291 5414 11343 5466
rect 11355 5414 11407 5466
rect 31526 5414 31578 5466
rect 31590 5414 31642 5466
rect 31654 5414 31706 5466
rect 31718 5414 31770 5466
rect 51888 5414 51940 5466
rect 51952 5414 52004 5466
rect 52016 5414 52068 5466
rect 52080 5414 52132 5466
rect 2964 5312 3016 5364
rect 6368 5312 6420 5364
rect 7012 5312 7064 5364
rect 12532 5355 12584 5364
rect 12532 5321 12541 5355
rect 12541 5321 12575 5355
rect 12575 5321 12584 5355
rect 12532 5312 12584 5321
rect 8392 5176 8444 5228
rect 14924 5312 14976 5364
rect 16672 5312 16724 5364
rect 17960 5312 18012 5364
rect 20904 5312 20956 5364
rect 23112 5312 23164 5364
rect 25504 5312 25556 5364
rect 36728 5312 36780 5364
rect 38016 5312 38068 5364
rect 40868 5312 40920 5364
rect 40960 5312 41012 5364
rect 11060 5176 11112 5228
rect 12256 5176 12308 5228
rect 23572 5244 23624 5296
rect 26884 5287 26936 5296
rect 2872 5151 2924 5160
rect 2872 5117 2901 5151
rect 2901 5117 2924 5151
rect 4160 5151 4212 5160
rect 2872 5108 2924 5117
rect 4160 5117 4169 5151
rect 4169 5117 4203 5151
rect 4203 5117 4212 5151
rect 4160 5108 4212 5117
rect 5356 5108 5408 5160
rect 7288 5108 7340 5160
rect 7840 5151 7892 5160
rect 7840 5117 7849 5151
rect 7849 5117 7883 5151
rect 7883 5117 7892 5151
rect 7840 5108 7892 5117
rect 8208 5108 8260 5160
rect 8944 5108 8996 5160
rect 9128 5108 9180 5160
rect 10876 5151 10928 5160
rect 10876 5117 10885 5151
rect 10885 5117 10919 5151
rect 10919 5117 10928 5151
rect 10876 5108 10928 5117
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 13728 5176 13780 5228
rect 15292 5219 15344 5228
rect 15292 5185 15301 5219
rect 15301 5185 15335 5219
rect 15335 5185 15344 5219
rect 15292 5176 15344 5185
rect 13544 5151 13596 5160
rect 13544 5117 13553 5151
rect 13553 5117 13587 5151
rect 13587 5117 13596 5151
rect 13544 5108 13596 5117
rect 5724 5040 5776 5092
rect 7932 4972 7984 5024
rect 14096 5040 14148 5092
rect 13728 4972 13780 5024
rect 15200 5108 15252 5160
rect 15752 5108 15804 5160
rect 16672 5151 16724 5160
rect 16672 5117 16681 5151
rect 16681 5117 16715 5151
rect 16715 5117 16724 5151
rect 16672 5108 16724 5117
rect 17224 5108 17276 5160
rect 20076 5219 20128 5228
rect 20076 5185 20085 5219
rect 20085 5185 20119 5219
rect 20119 5185 20128 5219
rect 20076 5176 20128 5185
rect 20628 5176 20680 5228
rect 26884 5253 26893 5287
rect 26893 5253 26927 5287
rect 26927 5253 26936 5287
rect 26884 5244 26936 5253
rect 26976 5244 27028 5296
rect 28448 5244 28500 5296
rect 24308 5176 24360 5228
rect 19892 5151 19944 5160
rect 18236 5083 18288 5092
rect 18236 5049 18245 5083
rect 18245 5049 18279 5083
rect 18279 5049 18288 5083
rect 18236 5040 18288 5049
rect 19892 5117 19901 5151
rect 19901 5117 19935 5151
rect 19935 5117 19944 5151
rect 19892 5108 19944 5117
rect 19984 5108 20036 5160
rect 24032 5151 24084 5160
rect 24032 5117 24041 5151
rect 24041 5117 24075 5151
rect 24075 5117 24084 5151
rect 24032 5108 24084 5117
rect 21180 5083 21232 5092
rect 15568 4972 15620 5024
rect 15660 4972 15712 5024
rect 17868 4972 17920 5024
rect 21180 5049 21189 5083
rect 21189 5049 21223 5083
rect 21223 5049 21232 5083
rect 21180 5040 21232 5049
rect 23664 5040 23716 5092
rect 25320 5108 25372 5160
rect 25504 5151 25556 5160
rect 25504 5117 25513 5151
rect 25513 5117 25547 5151
rect 25547 5117 25556 5151
rect 25504 5108 25556 5117
rect 25964 5151 26016 5160
rect 25964 5117 25973 5151
rect 25973 5117 26007 5151
rect 26007 5117 26016 5151
rect 25964 5108 26016 5117
rect 26608 5108 26660 5160
rect 32680 5176 32732 5228
rect 40592 5176 40644 5228
rect 40960 5176 41012 5228
rect 27712 5040 27764 5092
rect 31944 5151 31996 5160
rect 31944 5117 31953 5151
rect 31953 5117 31987 5151
rect 31987 5117 31996 5151
rect 32220 5151 32272 5160
rect 31944 5108 31996 5117
rect 32220 5117 32229 5151
rect 32229 5117 32263 5151
rect 32263 5117 32272 5151
rect 32220 5108 32272 5117
rect 32312 5108 32364 5160
rect 32496 5108 32548 5160
rect 33324 5151 33376 5160
rect 33324 5117 33333 5151
rect 33333 5117 33367 5151
rect 33367 5117 33376 5151
rect 33324 5108 33376 5117
rect 34796 5108 34848 5160
rect 36452 5151 36504 5160
rect 36452 5117 36461 5151
rect 36461 5117 36495 5151
rect 36495 5117 36504 5151
rect 36452 5108 36504 5117
rect 36544 5151 36596 5160
rect 36544 5117 36553 5151
rect 36553 5117 36587 5151
rect 36587 5117 36596 5151
rect 36728 5151 36780 5160
rect 36544 5108 36596 5117
rect 36728 5117 36737 5151
rect 36737 5117 36771 5151
rect 36771 5117 36780 5151
rect 36728 5108 36780 5117
rect 36912 5151 36964 5160
rect 36912 5117 36921 5151
rect 36921 5117 36955 5151
rect 36955 5117 36964 5151
rect 36912 5108 36964 5117
rect 37096 5108 37148 5160
rect 37188 5108 37240 5160
rect 39028 5151 39080 5160
rect 39028 5117 39037 5151
rect 39037 5117 39071 5151
rect 39071 5117 39080 5151
rect 39028 5108 39080 5117
rect 39120 5108 39172 5160
rect 39488 5108 39540 5160
rect 39672 5108 39724 5160
rect 40316 5108 40368 5160
rect 41604 5176 41656 5228
rect 41420 5151 41472 5160
rect 41420 5117 41429 5151
rect 41429 5117 41463 5151
rect 41463 5117 41472 5151
rect 41420 5108 41472 5117
rect 42248 5151 42300 5160
rect 42248 5117 42257 5151
rect 42257 5117 42291 5151
rect 42291 5117 42300 5151
rect 42248 5108 42300 5117
rect 32864 5040 32916 5092
rect 25964 4972 26016 5024
rect 28724 4972 28776 5024
rect 30564 4972 30616 5024
rect 38936 5040 38988 5092
rect 33416 4972 33468 5024
rect 34244 4972 34296 5024
rect 34888 4972 34940 5024
rect 36176 4972 36228 5024
rect 36912 4972 36964 5024
rect 51448 5312 51500 5364
rect 51540 5312 51592 5364
rect 53012 5355 53064 5364
rect 53012 5321 53021 5355
rect 53021 5321 53055 5355
rect 53055 5321 53064 5355
rect 53012 5312 53064 5321
rect 55312 5312 55364 5364
rect 57520 5312 57572 5364
rect 47676 5287 47728 5296
rect 47676 5253 47685 5287
rect 47685 5253 47719 5287
rect 47719 5253 47728 5287
rect 47676 5244 47728 5253
rect 50068 5287 50120 5296
rect 50068 5253 50077 5287
rect 50077 5253 50111 5287
rect 50111 5253 50120 5287
rect 50068 5244 50120 5253
rect 53472 5244 53524 5296
rect 45468 5176 45520 5228
rect 46388 5219 46440 5228
rect 46388 5185 46397 5219
rect 46397 5185 46431 5219
rect 46431 5185 46440 5219
rect 46388 5176 46440 5185
rect 43720 5151 43772 5160
rect 43720 5117 43729 5151
rect 43729 5117 43763 5151
rect 43763 5117 43772 5151
rect 43720 5108 43772 5117
rect 46112 5151 46164 5160
rect 46112 5117 46121 5151
rect 46121 5117 46155 5151
rect 46155 5117 46164 5151
rect 46112 5108 46164 5117
rect 46204 5108 46256 5160
rect 49608 5108 49660 5160
rect 49792 5151 49844 5160
rect 49792 5117 49801 5151
rect 49801 5117 49835 5151
rect 49835 5117 49844 5151
rect 49792 5108 49844 5117
rect 44180 5040 44232 5092
rect 47952 5040 48004 5092
rect 50436 5040 50488 5092
rect 49976 4972 50028 5024
rect 50528 4972 50580 5024
rect 50804 5176 50856 5228
rect 53380 5176 53432 5228
rect 53748 5108 53800 5160
rect 50712 5040 50764 5092
rect 54852 5108 54904 5160
rect 57980 5176 58032 5228
rect 58072 5176 58124 5228
rect 56508 5108 56560 5160
rect 55404 5083 55456 5092
rect 55404 5049 55413 5083
rect 55413 5049 55447 5083
rect 55447 5049 55456 5083
rect 55404 5040 55456 5049
rect 58440 5108 58492 5160
rect 21344 4870 21396 4922
rect 21408 4870 21460 4922
rect 21472 4870 21524 4922
rect 21536 4870 21588 4922
rect 41707 4870 41759 4922
rect 41771 4870 41823 4922
rect 41835 4870 41887 4922
rect 41899 4870 41951 4922
rect 6368 4768 6420 4820
rect 15200 4768 15252 4820
rect 3240 4700 3292 4752
rect 5356 4743 5408 4752
rect 5356 4709 5365 4743
rect 5365 4709 5399 4743
rect 5399 4709 5408 4743
rect 5356 4700 5408 4709
rect 2688 4675 2740 4684
rect 2688 4641 2697 4675
rect 2697 4641 2731 4675
rect 2731 4641 2740 4675
rect 2688 4632 2740 4641
rect 4068 4675 4120 4684
rect 4068 4641 4077 4675
rect 4077 4641 4111 4675
rect 4111 4641 4120 4675
rect 4068 4632 4120 4641
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 6920 4632 6972 4684
rect 8392 4700 8444 4752
rect 12440 4700 12492 4752
rect 8116 4675 8168 4684
rect 8116 4641 8125 4675
rect 8125 4641 8159 4675
rect 8159 4641 8168 4675
rect 8116 4632 8168 4641
rect 12164 4632 12216 4684
rect 13636 4743 13688 4752
rect 13636 4709 13645 4743
rect 13645 4709 13679 4743
rect 13679 4709 13688 4743
rect 16212 4768 16264 4820
rect 16948 4768 17000 4820
rect 13636 4700 13688 4709
rect 25228 4768 25280 4820
rect 28172 4768 28224 4820
rect 29000 4768 29052 4820
rect 30840 4768 30892 4820
rect 31944 4768 31996 4820
rect 7104 4564 7156 4616
rect 7380 4607 7432 4616
rect 7380 4573 7389 4607
rect 7389 4573 7423 4607
rect 7423 4573 7432 4607
rect 7380 4564 7432 4573
rect 13176 4632 13228 4684
rect 12808 4564 12860 4616
rect 12440 4496 12492 4548
rect 4160 4471 4212 4480
rect 4160 4437 4169 4471
rect 4169 4437 4203 4471
rect 4203 4437 4212 4471
rect 4160 4428 4212 4437
rect 8668 4428 8720 4480
rect 11980 4471 12032 4480
rect 11980 4437 11989 4471
rect 11989 4437 12023 4471
rect 12023 4437 12032 4471
rect 11980 4428 12032 4437
rect 13728 4632 13780 4684
rect 23112 4700 23164 4752
rect 16304 4632 16356 4684
rect 20996 4632 21048 4684
rect 22468 4675 22520 4684
rect 14004 4607 14056 4616
rect 14004 4573 14013 4607
rect 14013 4573 14047 4607
rect 14047 4573 14056 4607
rect 14004 4564 14056 4573
rect 15384 4564 15436 4616
rect 16672 4564 16724 4616
rect 16856 4607 16908 4616
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 17868 4607 17920 4616
rect 15752 4496 15804 4548
rect 16028 4496 16080 4548
rect 17868 4573 17877 4607
rect 17877 4573 17911 4607
rect 17911 4573 17920 4607
rect 17868 4564 17920 4573
rect 21916 4564 21968 4616
rect 22468 4641 22477 4675
rect 22477 4641 22511 4675
rect 22511 4641 22520 4675
rect 22468 4632 22520 4641
rect 22744 4675 22796 4684
rect 22744 4641 22753 4675
rect 22753 4641 22787 4675
rect 22787 4641 22796 4675
rect 22744 4632 22796 4641
rect 24860 4675 24912 4684
rect 22560 4564 22612 4616
rect 24308 4564 24360 4616
rect 18236 4496 18288 4548
rect 19248 4496 19300 4548
rect 24032 4496 24084 4548
rect 24860 4641 24869 4675
rect 24869 4641 24903 4675
rect 24903 4641 24912 4675
rect 24860 4632 24912 4641
rect 25412 4632 25464 4684
rect 26424 4632 26476 4684
rect 26976 4700 27028 4752
rect 29092 4700 29144 4752
rect 31116 4700 31168 4752
rect 29184 4632 29236 4684
rect 29736 4632 29788 4684
rect 31024 4675 31076 4684
rect 31024 4641 31033 4675
rect 31033 4641 31067 4675
rect 31067 4641 31076 4675
rect 31024 4632 31076 4641
rect 31944 4632 31996 4684
rect 32036 4632 32088 4684
rect 33140 4768 33192 4820
rect 43720 4768 43772 4820
rect 45744 4768 45796 4820
rect 32496 4632 32548 4684
rect 37188 4700 37240 4752
rect 38108 4700 38160 4752
rect 28632 4607 28684 4616
rect 28632 4573 28641 4607
rect 28641 4573 28675 4607
rect 28675 4573 28684 4607
rect 28632 4564 28684 4573
rect 30564 4564 30616 4616
rect 28908 4496 28960 4548
rect 36084 4564 36136 4616
rect 36360 4632 36412 4684
rect 38384 4675 38436 4684
rect 38384 4641 38393 4675
rect 38393 4641 38427 4675
rect 38427 4641 38436 4675
rect 38384 4632 38436 4641
rect 40040 4700 40092 4752
rect 38936 4632 38988 4684
rect 41972 4632 42024 4684
rect 35348 4539 35400 4548
rect 35348 4505 35357 4539
rect 35357 4505 35391 4539
rect 35391 4505 35400 4539
rect 35348 4496 35400 4505
rect 37280 4564 37332 4616
rect 40868 4564 40920 4616
rect 41236 4564 41288 4616
rect 37832 4496 37884 4548
rect 40408 4496 40460 4548
rect 45468 4632 45520 4684
rect 46572 4675 46624 4684
rect 46572 4641 46581 4675
rect 46581 4641 46615 4675
rect 46615 4641 46624 4675
rect 46572 4632 46624 4641
rect 47952 4743 48004 4752
rect 47952 4709 47961 4743
rect 47961 4709 47995 4743
rect 47995 4709 48004 4743
rect 50436 4768 50488 4820
rect 47952 4700 48004 4709
rect 50804 4700 50856 4752
rect 49056 4632 49108 4684
rect 51724 4632 51776 4684
rect 58624 4768 58676 4820
rect 58808 4768 58860 4820
rect 57612 4700 57664 4752
rect 52460 4675 52512 4684
rect 52460 4641 52469 4675
rect 52469 4641 52503 4675
rect 52503 4641 52512 4675
rect 52460 4632 52512 4641
rect 56324 4632 56376 4684
rect 56508 4675 56560 4684
rect 56508 4641 56517 4675
rect 56517 4641 56551 4675
rect 56551 4641 56560 4675
rect 60188 4700 60240 4752
rect 58808 4675 58860 4684
rect 56508 4632 56560 4641
rect 58808 4641 58817 4675
rect 58817 4641 58851 4675
rect 58851 4641 58860 4675
rect 58808 4632 58860 4641
rect 48780 4564 48832 4616
rect 49424 4564 49476 4616
rect 50436 4564 50488 4616
rect 52276 4564 52328 4616
rect 57980 4607 58032 4616
rect 55404 4496 55456 4548
rect 57980 4573 57989 4607
rect 57989 4573 58023 4607
rect 58023 4573 58032 4607
rect 57980 4564 58032 4573
rect 56692 4496 56744 4548
rect 58440 4539 58492 4548
rect 58440 4505 58449 4539
rect 58449 4505 58483 4539
rect 58483 4505 58492 4539
rect 58440 4496 58492 4505
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 18880 4428 18932 4480
rect 18972 4428 19024 4480
rect 20352 4428 20404 4480
rect 28356 4428 28408 4480
rect 28724 4428 28776 4480
rect 31024 4428 31076 4480
rect 31300 4428 31352 4480
rect 32036 4428 32088 4480
rect 33324 4428 33376 4480
rect 34980 4428 35032 4480
rect 37464 4428 37516 4480
rect 38108 4428 38160 4480
rect 38660 4471 38712 4480
rect 38660 4437 38669 4471
rect 38669 4437 38703 4471
rect 38703 4437 38712 4471
rect 38660 4428 38712 4437
rect 46940 4428 46992 4480
rect 55680 4428 55732 4480
rect 11163 4326 11215 4378
rect 11227 4326 11279 4378
rect 11291 4326 11343 4378
rect 11355 4326 11407 4378
rect 31526 4326 31578 4378
rect 31590 4326 31642 4378
rect 31654 4326 31706 4378
rect 31718 4326 31770 4378
rect 51888 4326 51940 4378
rect 51952 4326 52004 4378
rect 52016 4326 52068 4378
rect 52080 4326 52132 4378
rect 6920 4224 6972 4276
rect 8024 4224 8076 4276
rect 11980 4224 12032 4276
rect 13636 4224 13688 4276
rect 14004 4224 14056 4276
rect 22468 4224 22520 4276
rect 27804 4224 27856 4276
rect 28908 4224 28960 4276
rect 31392 4224 31444 4276
rect 32220 4224 32272 4276
rect 33048 4224 33100 4276
rect 37372 4224 37424 4276
rect 41052 4224 41104 4276
rect 46848 4224 46900 4276
rect 49700 4224 49752 4276
rect 51356 4224 51408 4276
rect 52276 4224 52328 4276
rect 6828 4156 6880 4208
rect 4528 4131 4580 4140
rect 2688 4063 2740 4072
rect 2688 4029 2697 4063
rect 2697 4029 2731 4063
rect 2731 4029 2740 4063
rect 3976 4063 4028 4072
rect 2688 4020 2740 4029
rect 3976 4029 3985 4063
rect 3985 4029 4019 4063
rect 4019 4029 4028 4063
rect 3976 4020 4028 4029
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 4528 4088 4580 4097
rect 7196 4088 7248 4140
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 9036 4088 9088 4140
rect 11060 4156 11112 4208
rect 11612 4156 11664 4208
rect 19984 4156 20036 4208
rect 13544 4088 13596 4140
rect 5356 4063 5408 4072
rect 5356 4029 5365 4063
rect 5365 4029 5399 4063
rect 5399 4029 5408 4063
rect 5356 4020 5408 4029
rect 5724 4020 5776 4072
rect 7472 4063 7524 4072
rect 7472 4029 7481 4063
rect 7481 4029 7515 4063
rect 7515 4029 7524 4063
rect 7472 4020 7524 4029
rect 7564 3952 7616 4004
rect 6736 3884 6788 3936
rect 6920 3927 6972 3936
rect 6920 3893 6929 3927
rect 6929 3893 6963 3927
rect 6963 3893 6972 3927
rect 6920 3884 6972 3893
rect 8668 3952 8720 4004
rect 9956 3952 10008 4004
rect 13176 4063 13228 4072
rect 13176 4029 13185 4063
rect 13185 4029 13219 4063
rect 13219 4029 13228 4063
rect 15200 4088 15252 4140
rect 18236 4131 18288 4140
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 20168 4131 20220 4140
rect 20168 4097 20177 4131
rect 20177 4097 20211 4131
rect 20211 4097 20220 4131
rect 20168 4088 20220 4097
rect 22560 4088 22612 4140
rect 24860 4088 24912 4140
rect 13176 4020 13228 4029
rect 13268 3952 13320 4004
rect 14188 4020 14240 4072
rect 15292 4063 15344 4072
rect 15292 4029 15301 4063
rect 15301 4029 15335 4063
rect 15335 4029 15344 4063
rect 15292 4020 15344 4029
rect 16672 4063 16724 4072
rect 16672 4029 16681 4063
rect 16681 4029 16715 4063
rect 16715 4029 16724 4063
rect 16672 4020 16724 4029
rect 16856 4020 16908 4072
rect 17224 4020 17276 4072
rect 18788 4020 18840 4072
rect 19064 4063 19116 4072
rect 19064 4029 19095 4063
rect 19095 4029 19116 4063
rect 19064 4020 19116 4029
rect 19248 4020 19300 4072
rect 20076 4063 20128 4072
rect 20076 4029 20085 4063
rect 20085 4029 20119 4063
rect 20119 4029 20128 4063
rect 20076 4020 20128 4029
rect 20352 4063 20404 4072
rect 20352 4029 20361 4063
rect 20361 4029 20395 4063
rect 20395 4029 20404 4063
rect 20352 4020 20404 4029
rect 13452 3952 13504 4004
rect 16028 3952 16080 4004
rect 18328 3995 18380 4004
rect 9128 3884 9180 3936
rect 18328 3961 18337 3995
rect 18337 3961 18371 3995
rect 18371 3961 18380 3995
rect 18328 3952 18380 3961
rect 23664 4020 23716 4072
rect 23848 4063 23900 4072
rect 23848 4029 23857 4063
rect 23857 4029 23891 4063
rect 23891 4029 23900 4063
rect 28264 4088 28316 4140
rect 34980 4156 35032 4208
rect 37740 4156 37792 4208
rect 31208 4088 31260 4140
rect 23848 4020 23900 4029
rect 26056 4020 26108 4072
rect 20812 3952 20864 4004
rect 23296 3952 23348 4004
rect 26792 3952 26844 4004
rect 29000 4020 29052 4072
rect 29276 4020 29328 4072
rect 29552 4020 29604 4072
rect 31024 4020 31076 4072
rect 31300 4020 31352 4072
rect 30104 3995 30156 4004
rect 30104 3961 30113 3995
rect 30113 3961 30147 3995
rect 30147 3961 30156 3995
rect 30104 3952 30156 3961
rect 30932 3952 30984 4004
rect 31116 3952 31168 4004
rect 34980 4020 35032 4072
rect 36084 4020 36136 4072
rect 37280 4063 37332 4072
rect 32496 3952 32548 4004
rect 37280 4029 37289 4063
rect 37289 4029 37323 4063
rect 37323 4029 37332 4063
rect 37280 4020 37332 4029
rect 37464 4088 37516 4140
rect 37924 4088 37976 4140
rect 38568 4088 38620 4140
rect 38936 4088 38988 4140
rect 40040 4088 40092 4140
rect 45744 4156 45796 4208
rect 49424 4199 49476 4208
rect 40500 4088 40552 4140
rect 40868 4131 40920 4140
rect 40868 4097 40877 4131
rect 40877 4097 40911 4131
rect 40911 4097 40920 4131
rect 40868 4088 40920 4097
rect 45560 4088 45612 4140
rect 49424 4165 49433 4199
rect 49433 4165 49467 4199
rect 49467 4165 49476 4199
rect 49424 4156 49476 4165
rect 39304 4020 39356 4072
rect 39580 4063 39632 4072
rect 39580 4029 39589 4063
rect 39589 4029 39623 4063
rect 39623 4029 39632 4063
rect 39580 4020 39632 4029
rect 43076 4020 43128 4072
rect 44916 4063 44968 4072
rect 36636 3952 36688 4004
rect 38200 3952 38252 4004
rect 39212 3952 39264 4004
rect 44916 4029 44925 4063
rect 44925 4029 44959 4063
rect 44959 4029 44968 4063
rect 44916 4020 44968 4029
rect 45468 4020 45520 4072
rect 18788 3884 18840 3936
rect 18880 3884 18932 3936
rect 20076 3884 20128 3936
rect 20536 3927 20588 3936
rect 20536 3893 20545 3927
rect 20545 3893 20579 3927
rect 20579 3893 20588 3927
rect 20536 3884 20588 3893
rect 22652 3927 22704 3936
rect 22652 3893 22661 3927
rect 22661 3893 22695 3927
rect 22695 3893 22704 3927
rect 22652 3884 22704 3893
rect 27252 3927 27304 3936
rect 27252 3893 27261 3927
rect 27261 3893 27295 3927
rect 27295 3893 27304 3927
rect 27252 3884 27304 3893
rect 27344 3884 27396 3936
rect 31852 3884 31904 3936
rect 32036 3884 32088 3936
rect 32680 3884 32732 3936
rect 34428 3884 34480 3936
rect 35716 3884 35768 3936
rect 36176 3884 36228 3936
rect 41144 3884 41196 3936
rect 41236 3884 41288 3936
rect 46572 3952 46624 4004
rect 47584 4020 47636 4072
rect 49516 4020 49568 4072
rect 51724 4088 51776 4140
rect 49884 4020 49936 4072
rect 50068 4020 50120 4072
rect 48228 3952 48280 4004
rect 54024 4088 54076 4140
rect 55312 4088 55364 4140
rect 56692 4088 56744 4140
rect 53472 4020 53524 4072
rect 55404 4063 55456 4072
rect 55404 4029 55413 4063
rect 55413 4029 55447 4063
rect 55447 4029 55456 4063
rect 55404 4020 55456 4029
rect 55864 4063 55916 4072
rect 55864 4029 55873 4063
rect 55873 4029 55907 4063
rect 55907 4029 55916 4063
rect 55864 4020 55916 4029
rect 55956 4020 56008 4072
rect 59452 4088 59504 4140
rect 57796 4020 57848 4072
rect 58532 4063 58584 4072
rect 58532 4029 58541 4063
rect 58541 4029 58575 4063
rect 58575 4029 58584 4063
rect 58532 4020 58584 4029
rect 58808 4063 58860 4072
rect 58808 4029 58817 4063
rect 58817 4029 58851 4063
rect 58851 4029 58860 4063
rect 58808 4020 58860 4029
rect 45652 3884 45704 3936
rect 51632 3884 51684 3936
rect 53748 3884 53800 3936
rect 55588 3884 55640 3936
rect 55956 3884 56008 3936
rect 57704 3884 57756 3936
rect 57980 3884 58032 3936
rect 21344 3782 21396 3834
rect 21408 3782 21460 3834
rect 21472 3782 21524 3834
rect 21536 3782 21588 3834
rect 41707 3782 41759 3834
rect 41771 3782 41823 3834
rect 41835 3782 41887 3834
rect 41899 3782 41951 3834
rect 3976 3680 4028 3732
rect 14188 3680 14240 3732
rect 16028 3680 16080 3732
rect 19064 3680 19116 3732
rect 21088 3723 21140 3732
rect 21088 3689 21097 3723
rect 21097 3689 21131 3723
rect 21131 3689 21140 3723
rect 21088 3680 21140 3689
rect 23480 3723 23532 3732
rect 23480 3689 23489 3723
rect 23489 3689 23523 3723
rect 23523 3689 23532 3723
rect 23480 3680 23532 3689
rect 25504 3680 25556 3732
rect 27344 3680 27396 3732
rect 27804 3723 27856 3732
rect 27804 3689 27813 3723
rect 27813 3689 27847 3723
rect 27847 3689 27856 3723
rect 27804 3680 27856 3689
rect 6644 3612 6696 3664
rect 6736 3612 6788 3664
rect 12716 3612 12768 3664
rect 12992 3612 13044 3664
rect 22652 3612 22704 3664
rect 27712 3655 27764 3664
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 4988 3519 5040 3528
rect 4988 3485 4997 3519
rect 4997 3485 5031 3519
rect 5031 3485 5040 3519
rect 4988 3476 5040 3485
rect 6552 3519 6604 3528
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 7380 3544 7432 3596
rect 7932 3587 7984 3596
rect 7932 3553 7941 3587
rect 7941 3553 7975 3587
rect 7975 3553 7984 3587
rect 7932 3544 7984 3553
rect 8576 3587 8628 3596
rect 8576 3553 8585 3587
rect 8585 3553 8619 3587
rect 8619 3553 8628 3587
rect 8576 3544 8628 3553
rect 12808 3544 12860 3596
rect 13084 3587 13136 3596
rect 13084 3553 13093 3587
rect 13093 3553 13127 3587
rect 13127 3553 13136 3587
rect 13084 3544 13136 3553
rect 16304 3587 16356 3596
rect 8208 3476 8260 3528
rect 10784 3476 10836 3528
rect 12440 3476 12492 3528
rect 16304 3553 16313 3587
rect 16313 3553 16347 3587
rect 16347 3553 16356 3587
rect 16304 3544 16356 3553
rect 13728 3476 13780 3528
rect 15568 3476 15620 3528
rect 16856 3544 16908 3596
rect 17224 3587 17276 3596
rect 17224 3553 17233 3587
rect 17233 3553 17267 3587
rect 17267 3553 17276 3587
rect 18880 3587 18932 3596
rect 17224 3544 17276 3553
rect 17500 3476 17552 3528
rect 18512 3476 18564 3528
rect 5356 3408 5408 3460
rect 5540 3340 5592 3392
rect 7472 3408 7524 3460
rect 7840 3408 7892 3460
rect 8024 3408 8076 3460
rect 16028 3408 16080 3460
rect 16304 3408 16356 3460
rect 17776 3408 17828 3460
rect 18236 3408 18288 3460
rect 18880 3553 18889 3587
rect 18889 3553 18923 3587
rect 18923 3553 18932 3587
rect 18880 3544 18932 3553
rect 19248 3544 19300 3596
rect 19340 3587 19392 3596
rect 19340 3553 19349 3587
rect 19349 3553 19383 3587
rect 19383 3553 19392 3587
rect 20904 3587 20956 3596
rect 19340 3544 19392 3553
rect 20904 3553 20913 3587
rect 20913 3553 20947 3587
rect 20947 3553 20956 3587
rect 20904 3544 20956 3553
rect 23204 3587 23256 3596
rect 23204 3553 23213 3587
rect 23213 3553 23247 3587
rect 23247 3553 23256 3587
rect 23204 3544 23256 3553
rect 20720 3476 20772 3528
rect 22836 3476 22888 3528
rect 24216 3544 24268 3596
rect 27712 3621 27721 3655
rect 27721 3621 27755 3655
rect 27755 3621 27764 3655
rect 27712 3612 27764 3621
rect 27896 3655 27948 3664
rect 27896 3621 27905 3655
rect 27905 3621 27939 3655
rect 27939 3621 27948 3655
rect 27896 3612 27948 3621
rect 28264 3655 28316 3664
rect 28264 3621 28273 3655
rect 28273 3621 28307 3655
rect 28307 3621 28316 3655
rect 28264 3612 28316 3621
rect 24860 3476 24912 3528
rect 9128 3340 9180 3392
rect 13268 3340 13320 3392
rect 13912 3340 13964 3392
rect 20628 3408 20680 3460
rect 26240 3476 26292 3528
rect 27528 3519 27580 3528
rect 27528 3485 27537 3519
rect 27537 3485 27571 3519
rect 27571 3485 27580 3519
rect 27528 3476 27580 3485
rect 29736 3612 29788 3664
rect 30104 3680 30156 3732
rect 30012 3544 30064 3596
rect 31116 3476 31168 3528
rect 32312 3476 32364 3528
rect 39580 3680 39632 3732
rect 41604 3723 41656 3732
rect 41604 3689 41613 3723
rect 41613 3689 41647 3723
rect 41647 3689 41656 3723
rect 41604 3680 41656 3689
rect 43352 3680 43404 3732
rect 49700 3680 49752 3732
rect 49884 3723 49936 3732
rect 49884 3689 49893 3723
rect 49893 3689 49927 3723
rect 49927 3689 49936 3723
rect 49884 3680 49936 3689
rect 57612 3680 57664 3732
rect 33048 3519 33100 3528
rect 33048 3485 33057 3519
rect 33057 3485 33091 3519
rect 33091 3485 33100 3519
rect 34612 3612 34664 3664
rect 34428 3587 34480 3596
rect 33048 3476 33100 3485
rect 30564 3408 30616 3460
rect 30748 3408 30800 3460
rect 19708 3340 19760 3392
rect 20352 3340 20404 3392
rect 22468 3340 22520 3392
rect 29276 3340 29328 3392
rect 29368 3340 29420 3392
rect 31300 3340 31352 3392
rect 32404 3340 32456 3392
rect 32956 3340 33008 3392
rect 34428 3553 34437 3587
rect 34437 3553 34471 3587
rect 34471 3553 34480 3587
rect 34428 3544 34480 3553
rect 36176 3612 36228 3664
rect 36268 3612 36320 3664
rect 38844 3612 38896 3664
rect 55864 3612 55916 3664
rect 58808 3612 58860 3664
rect 35532 3519 35584 3528
rect 35532 3485 35541 3519
rect 35541 3485 35575 3519
rect 35575 3485 35584 3519
rect 35532 3476 35584 3485
rect 36360 3476 36412 3528
rect 36728 3544 36780 3596
rect 37188 3544 37240 3596
rect 37832 3544 37884 3596
rect 39028 3544 39080 3596
rect 39212 3587 39264 3596
rect 39212 3553 39221 3587
rect 39221 3553 39255 3587
rect 39255 3553 39264 3587
rect 39212 3544 39264 3553
rect 40408 3544 40460 3596
rect 43628 3544 43680 3596
rect 44088 3544 44140 3596
rect 46572 3587 46624 3596
rect 46572 3553 46581 3587
rect 46581 3553 46615 3587
rect 46615 3553 46624 3587
rect 46572 3544 46624 3553
rect 38476 3476 38528 3528
rect 37648 3340 37700 3392
rect 38568 3408 38620 3460
rect 40500 3476 40552 3528
rect 46112 3476 46164 3528
rect 49700 3544 49752 3596
rect 51632 3587 51684 3596
rect 51632 3553 51641 3587
rect 51641 3553 51675 3587
rect 51675 3553 51684 3587
rect 51632 3544 51684 3553
rect 55312 3587 55364 3596
rect 55312 3553 55321 3587
rect 55321 3553 55355 3587
rect 55355 3553 55364 3587
rect 55312 3544 55364 3553
rect 55680 3587 55732 3596
rect 55680 3553 55689 3587
rect 55689 3553 55723 3587
rect 55723 3553 55732 3587
rect 55680 3544 55732 3553
rect 56784 3587 56836 3596
rect 56784 3553 56793 3587
rect 56793 3553 56827 3587
rect 56827 3553 56836 3587
rect 56784 3544 56836 3553
rect 56876 3544 56928 3596
rect 58716 3587 58768 3596
rect 58716 3553 58725 3587
rect 58725 3553 58759 3587
rect 58759 3553 58768 3587
rect 58716 3544 58768 3553
rect 58900 3544 58952 3596
rect 61016 3544 61068 3596
rect 50436 3476 50488 3528
rect 51264 3476 51316 3528
rect 52184 3476 52236 3528
rect 53196 3476 53248 3528
rect 41144 3408 41196 3460
rect 43812 3408 43864 3460
rect 50620 3408 50672 3460
rect 54576 3476 54628 3528
rect 55588 3519 55640 3528
rect 55588 3485 55597 3519
rect 55597 3485 55631 3519
rect 55631 3485 55640 3519
rect 55588 3476 55640 3485
rect 55772 3476 55824 3528
rect 58440 3476 58492 3528
rect 41236 3340 41288 3392
rect 49976 3340 50028 3392
rect 51540 3340 51592 3392
rect 53564 3383 53616 3392
rect 53564 3349 53573 3383
rect 53573 3349 53607 3383
rect 53607 3349 53616 3383
rect 53564 3340 53616 3349
rect 58716 3340 58768 3392
rect 11163 3238 11215 3290
rect 11227 3238 11279 3290
rect 11291 3238 11343 3290
rect 11355 3238 11407 3290
rect 31526 3238 31578 3290
rect 31590 3238 31642 3290
rect 31654 3238 31706 3290
rect 31718 3238 31770 3290
rect 51888 3238 51940 3290
rect 51952 3238 52004 3290
rect 52016 3238 52068 3290
rect 52080 3238 52132 3290
rect 6460 3136 6512 3188
rect 4988 3000 5040 3052
rect 6552 3068 6604 3120
rect 7564 3136 7616 3188
rect 12992 3136 13044 3188
rect 13084 3136 13136 3188
rect 6920 3000 6972 3052
rect 7840 3043 7892 3052
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 8208 3000 8260 3052
rect 9864 3000 9916 3052
rect 13176 3068 13228 3120
rect 17592 3068 17644 3120
rect 17776 3136 17828 3188
rect 21180 3136 21232 3188
rect 22468 3136 22520 3188
rect 23664 3136 23716 3188
rect 26056 3136 26108 3188
rect 28080 3136 28132 3188
rect 33232 3136 33284 3188
rect 33324 3136 33376 3188
rect 5908 2864 5960 2916
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 8024 2932 8076 2984
rect 8116 2932 8168 2984
rect 13452 3043 13504 3052
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 12900 2864 12952 2916
rect 13728 2975 13780 2984
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 13912 2975 13964 2984
rect 13728 2932 13780 2941
rect 13912 2941 13921 2975
rect 13921 2941 13955 2975
rect 13955 2941 13964 2975
rect 13912 2932 13964 2941
rect 14740 2975 14792 2984
rect 14740 2941 14749 2975
rect 14749 2941 14783 2975
rect 14783 2941 14792 2975
rect 14740 2932 14792 2941
rect 16764 2932 16816 2984
rect 7288 2796 7340 2848
rect 16304 2796 16356 2848
rect 16580 2796 16632 2848
rect 18236 3000 18288 3052
rect 18328 3000 18380 3052
rect 24124 3068 24176 3120
rect 27528 3068 27580 3120
rect 21824 3000 21876 3052
rect 24860 3043 24912 3052
rect 24860 3009 24869 3043
rect 24869 3009 24903 3043
rect 24903 3009 24912 3043
rect 24860 3000 24912 3009
rect 16948 2975 17000 2984
rect 16948 2941 16957 2975
rect 16957 2941 16991 2975
rect 16991 2941 17000 2975
rect 16948 2932 17000 2941
rect 18696 2975 18748 2984
rect 17316 2864 17368 2916
rect 18696 2941 18705 2975
rect 18705 2941 18739 2975
rect 18739 2941 18748 2975
rect 18696 2932 18748 2941
rect 18788 2975 18840 2984
rect 18788 2941 18797 2975
rect 18797 2941 18831 2975
rect 18831 2941 18840 2975
rect 19064 2975 19116 2984
rect 18788 2932 18840 2941
rect 19064 2941 19073 2975
rect 19073 2941 19107 2975
rect 19107 2941 19116 2975
rect 19064 2932 19116 2941
rect 19248 2932 19300 2984
rect 20628 2932 20680 2984
rect 20812 2932 20864 2984
rect 22560 2932 22612 2984
rect 24308 2932 24360 2984
rect 34888 3068 34940 3120
rect 35992 3068 36044 3120
rect 28356 3043 28408 3052
rect 28356 3009 28365 3043
rect 28365 3009 28399 3043
rect 28399 3009 28408 3043
rect 28356 3000 28408 3009
rect 29000 3000 29052 3052
rect 30288 3000 30340 3052
rect 30472 3043 30524 3052
rect 30472 3009 30481 3043
rect 30481 3009 30515 3043
rect 30515 3009 30524 3043
rect 30472 3000 30524 3009
rect 30932 3043 30984 3052
rect 30932 3009 30941 3043
rect 30941 3009 30975 3043
rect 30975 3009 30984 3043
rect 30932 3000 30984 3009
rect 31024 3000 31076 3052
rect 32128 3000 32180 3052
rect 27896 2975 27948 2984
rect 27896 2941 27905 2975
rect 27905 2941 27939 2975
rect 27939 2941 27948 2975
rect 27896 2932 27948 2941
rect 30012 2932 30064 2984
rect 30748 2975 30800 2984
rect 30748 2941 30757 2975
rect 30757 2941 30791 2975
rect 30791 2941 30800 2975
rect 30748 2932 30800 2941
rect 26240 2907 26292 2916
rect 26240 2873 26249 2907
rect 26249 2873 26283 2907
rect 26283 2873 26292 2907
rect 26240 2864 26292 2873
rect 17960 2796 18012 2848
rect 18788 2796 18840 2848
rect 22836 2796 22888 2848
rect 30288 2864 30340 2916
rect 30380 2864 30432 2916
rect 32680 2932 32732 2984
rect 34336 3000 34388 3052
rect 34612 3000 34664 3052
rect 36636 3068 36688 3120
rect 36728 3000 36780 3052
rect 38108 3136 38160 3188
rect 38200 3043 38252 3052
rect 32956 2975 33008 2984
rect 32956 2941 32965 2975
rect 32965 2941 32999 2975
rect 32999 2941 33008 2975
rect 32956 2932 33008 2941
rect 35624 2932 35676 2984
rect 35716 2975 35768 2984
rect 35716 2941 35725 2975
rect 35725 2941 35759 2975
rect 35759 2941 35768 2975
rect 37924 2975 37976 2984
rect 35716 2932 35768 2941
rect 31392 2864 31444 2916
rect 36268 2864 36320 2916
rect 33048 2796 33100 2848
rect 35992 2839 36044 2848
rect 35992 2805 36001 2839
rect 36001 2805 36035 2839
rect 36035 2805 36044 2839
rect 37924 2941 37933 2975
rect 37933 2941 37967 2975
rect 37967 2941 37976 2975
rect 37924 2932 37976 2941
rect 38200 3009 38209 3043
rect 38209 3009 38243 3043
rect 38243 3009 38252 3043
rect 38200 3000 38252 3009
rect 39120 3000 39172 3052
rect 41512 3136 41564 3188
rect 40776 3111 40828 3120
rect 40776 3077 40785 3111
rect 40785 3077 40819 3111
rect 40819 3077 40828 3111
rect 40776 3068 40828 3077
rect 47032 3136 47084 3188
rect 38476 2932 38528 2984
rect 40500 2907 40552 2916
rect 40500 2873 40509 2907
rect 40509 2873 40543 2907
rect 40543 2873 40552 2907
rect 40500 2864 40552 2873
rect 41328 2932 41380 2984
rect 42064 2975 42116 2984
rect 42064 2941 42073 2975
rect 42073 2941 42107 2975
rect 42107 2941 42116 2975
rect 42064 2932 42116 2941
rect 45192 2932 45244 2984
rect 51264 3136 51316 3188
rect 52460 3179 52512 3188
rect 52460 3145 52469 3179
rect 52469 3145 52503 3179
rect 52503 3145 52512 3179
rect 52460 3136 52512 3145
rect 53472 3179 53524 3188
rect 53472 3145 53481 3179
rect 53481 3145 53515 3179
rect 53515 3145 53524 3179
rect 53472 3136 53524 3145
rect 53564 3136 53616 3188
rect 57980 3068 58032 3120
rect 61936 3068 61988 3120
rect 47032 2975 47084 2984
rect 44640 2907 44692 2916
rect 44640 2873 44649 2907
rect 44649 2873 44683 2907
rect 44683 2873 44692 2907
rect 44640 2864 44692 2873
rect 47032 2941 47041 2975
rect 47041 2941 47075 2975
rect 47075 2941 47084 2975
rect 47032 2932 47084 2941
rect 35992 2796 36044 2805
rect 43352 2796 43404 2848
rect 44088 2796 44140 2848
rect 52184 3000 52236 3052
rect 55404 3000 55456 3052
rect 58716 3043 58768 3052
rect 58716 3009 58725 3043
rect 58725 3009 58759 3043
rect 58759 3009 58768 3043
rect 58716 3000 58768 3009
rect 47584 2932 47636 2984
rect 49792 2932 49844 2984
rect 49976 2975 50028 2984
rect 49976 2941 49985 2975
rect 49985 2941 50019 2975
rect 50019 2941 50028 2975
rect 49976 2932 50028 2941
rect 53748 2932 53800 2984
rect 54024 2975 54076 2984
rect 54024 2941 54033 2975
rect 54033 2941 54067 2975
rect 54067 2941 54076 2975
rect 54024 2932 54076 2941
rect 54392 2975 54444 2984
rect 54392 2941 54401 2975
rect 54401 2941 54435 2975
rect 54435 2941 54444 2975
rect 54392 2932 54444 2941
rect 54576 2975 54628 2984
rect 54576 2941 54585 2975
rect 54585 2941 54619 2975
rect 54619 2941 54628 2975
rect 54576 2932 54628 2941
rect 54668 2932 54720 2984
rect 55588 2975 55640 2984
rect 55588 2941 55597 2975
rect 55597 2941 55631 2975
rect 55631 2941 55640 2975
rect 55588 2932 55640 2941
rect 56692 2932 56744 2984
rect 48504 2796 48556 2848
rect 49792 2796 49844 2848
rect 54668 2796 54720 2848
rect 56784 2864 56836 2916
rect 59268 2864 59320 2916
rect 60648 2796 60700 2848
rect 62764 2796 62816 2848
rect 21344 2694 21396 2746
rect 21408 2694 21460 2746
rect 21472 2694 21524 2746
rect 21536 2694 21588 2746
rect 41707 2694 41759 2746
rect 41771 2694 41823 2746
rect 41835 2694 41887 2746
rect 41899 2694 41951 2746
rect 2044 2456 2096 2508
rect 22100 2592 22152 2644
rect 30012 2592 30064 2644
rect 6828 2524 6880 2576
rect 8668 2524 8720 2576
rect 20812 2524 20864 2576
rect 26056 2524 26108 2576
rect 2964 2499 3016 2508
rect 2964 2465 2973 2499
rect 2973 2465 3007 2499
rect 3007 2465 3016 2499
rect 2964 2456 3016 2465
rect 5540 2456 5592 2508
rect 5908 2456 5960 2508
rect 12348 2456 12400 2508
rect 12900 2499 12952 2508
rect 12900 2465 12909 2499
rect 12909 2465 12943 2499
rect 12943 2465 12952 2499
rect 12900 2456 12952 2465
rect 17316 2456 17368 2508
rect 17592 2456 17644 2508
rect 21088 2456 21140 2508
rect 4344 2431 4396 2440
rect 4344 2397 4353 2431
rect 4353 2397 4387 2431
rect 4387 2397 4396 2431
rect 4344 2388 4396 2397
rect 12808 2388 12860 2440
rect 16396 2388 16448 2440
rect 16672 2388 16724 2440
rect 18328 2431 18380 2440
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18328 2388 18380 2397
rect 19708 2431 19760 2440
rect 19708 2397 19717 2431
rect 19717 2397 19751 2431
rect 19751 2397 19760 2431
rect 19708 2388 19760 2397
rect 20720 2388 20772 2440
rect 22836 2456 22888 2508
rect 26884 2499 26936 2508
rect 26884 2465 26893 2499
rect 26893 2465 26927 2499
rect 26927 2465 26936 2499
rect 26884 2456 26936 2465
rect 31024 2524 31076 2576
rect 32588 2524 32640 2576
rect 28264 2456 28316 2508
rect 30288 2499 30340 2508
rect 30288 2465 30297 2499
rect 30297 2465 30331 2499
rect 30331 2465 30340 2499
rect 30288 2456 30340 2465
rect 41512 2592 41564 2644
rect 44640 2592 44692 2644
rect 45192 2592 45244 2644
rect 48596 2592 48648 2644
rect 57980 2592 58032 2644
rect 33968 2567 34020 2576
rect 33968 2533 33977 2567
rect 33977 2533 34011 2567
rect 34011 2533 34020 2567
rect 33968 2524 34020 2533
rect 38108 2524 38160 2576
rect 40776 2524 40828 2576
rect 58440 2524 58492 2576
rect 35900 2499 35952 2508
rect 24308 2431 24360 2440
rect 24308 2397 24317 2431
rect 24317 2397 24351 2431
rect 24351 2397 24360 2431
rect 24308 2388 24360 2397
rect 17960 2252 18012 2304
rect 21732 2252 21784 2304
rect 24952 2252 25004 2304
rect 31116 2388 31168 2440
rect 32772 2388 32824 2440
rect 34612 2388 34664 2440
rect 35900 2465 35909 2499
rect 35909 2465 35943 2499
rect 35943 2465 35952 2499
rect 35900 2456 35952 2465
rect 36268 2499 36320 2508
rect 36268 2465 36277 2499
rect 36277 2465 36311 2499
rect 36311 2465 36320 2499
rect 36268 2456 36320 2465
rect 37924 2456 37976 2508
rect 38660 2456 38712 2508
rect 41052 2456 41104 2508
rect 41328 2456 41380 2508
rect 44548 2456 44600 2508
rect 48044 2456 48096 2508
rect 48504 2499 48556 2508
rect 48504 2465 48513 2499
rect 48513 2465 48547 2499
rect 48547 2465 48556 2499
rect 48504 2456 48556 2465
rect 54944 2456 54996 2508
rect 36084 2388 36136 2440
rect 40224 2388 40276 2440
rect 43720 2388 43772 2440
rect 47124 2388 47176 2440
rect 49792 2388 49844 2440
rect 60188 2456 60240 2508
rect 57612 2388 57664 2440
rect 41972 2320 42024 2372
rect 45468 2320 45520 2372
rect 46296 2320 46348 2372
rect 60648 2320 60700 2372
rect 29736 2252 29788 2304
rect 32864 2295 32916 2304
rect 32864 2261 32873 2295
rect 32873 2261 32907 2295
rect 32907 2261 32916 2295
rect 32864 2252 32916 2261
rect 39488 2252 39540 2304
rect 42800 2295 42852 2304
rect 42800 2261 42809 2295
rect 42809 2261 42843 2295
rect 42843 2261 42852 2295
rect 42800 2252 42852 2261
rect 42892 2252 42944 2304
rect 48872 2252 48924 2304
rect 52368 2252 52420 2304
rect 54116 2252 54168 2304
rect 11163 2150 11215 2202
rect 11227 2150 11279 2202
rect 11291 2150 11343 2202
rect 11355 2150 11407 2202
rect 31526 2150 31578 2202
rect 31590 2150 31642 2202
rect 31654 2150 31706 2202
rect 31718 2150 31770 2202
rect 51888 2150 51940 2202
rect 51952 2150 52004 2202
rect 52016 2150 52068 2202
rect 52080 2150 52132 2202
rect 16396 2048 16448 2100
rect 18328 2048 18380 2100
rect 21732 2048 21784 2100
rect 22100 2048 22152 2100
rect 31024 2048 31076 2100
rect 32588 2048 32640 2100
rect 40500 2048 40552 2100
rect 14464 1980 14516 2032
rect 16856 1980 16908 2032
rect 36268 1980 36320 2032
rect 37648 1980 37700 2032
rect 12716 1912 12768 1964
rect 13360 1912 13412 1964
rect 18972 1912 19024 1964
rect 36360 1912 36412 1964
rect 42800 1980 42852 2032
rect 32772 1844 32824 1896
rect 34796 1844 34848 1896
rect 38476 1844 38528 1896
rect 36084 1776 36136 1828
rect 36728 1776 36780 1828
rect 3424 1300 3476 1352
rect 27160 1300 27212 1352
<< metal2 >>
rect 938 18835 994 19635
rect 2778 18835 2834 19635
rect 4710 18835 4766 19635
rect 6642 18835 6698 19635
rect 8574 18835 8630 19635
rect 10506 18835 10562 19635
rect 12438 18835 12494 19635
rect 14278 18835 14334 19635
rect 16210 18835 16266 19635
rect 18142 18835 18198 19635
rect 20074 18835 20130 19635
rect 22006 18835 22062 19635
rect 23938 18835 23994 19635
rect 25870 18835 25926 19635
rect 27710 18835 27766 19635
rect 29642 18835 29698 19635
rect 31574 18835 31630 19635
rect 33506 18835 33562 19635
rect 35438 18835 35494 19635
rect 37370 18835 37426 19635
rect 39210 18835 39266 19635
rect 41142 18835 41198 19635
rect 43074 18835 43130 19635
rect 45006 18835 45062 19635
rect 46938 18835 46994 19635
rect 48870 18835 48926 19635
rect 50802 18835 50858 19635
rect 52642 18835 52698 19635
rect 54574 18835 54630 19635
rect 56506 18835 56562 19635
rect 58438 18835 58494 19635
rect 60370 18835 60426 19635
rect 62302 18835 62358 19635
rect 952 15910 980 18835
rect 2792 15978 2820 18835
rect 3330 18592 3386 18601
rect 3330 18527 3386 18536
rect 3054 16416 3110 16425
rect 3054 16351 3110 16360
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 940 15904 992 15910
rect 940 15846 992 15852
rect 3068 12918 3096 16351
rect 3344 13734 3372 18527
rect 4724 15638 4752 18835
rect 4712 15632 4764 15638
rect 4712 15574 4764 15580
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 4066 14240 4122 14249
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 3056 12912 3108 12918
rect 3056 12854 3108 12860
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2792 11218 2820 12378
rect 3528 12073 3556 14214
rect 4066 14175 4122 14184
rect 4080 13530 4108 14175
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5276 13870 5304 14010
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 5276 13394 5304 13806
rect 5368 13462 5396 15302
rect 5460 14958 5488 15438
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5460 12986 5488 13330
rect 5552 13190 5580 14350
rect 5644 13938 5672 14758
rect 6012 14618 6040 15506
rect 6656 14958 6684 18835
rect 8116 15632 8168 15638
rect 8116 15574 8168 15580
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 6656 14618 6684 14894
rect 6000 14612 6052 14618
rect 6000 14554 6052 14560
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 7024 13870 7052 15302
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7116 14482 7144 14894
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 14006 7328 14214
rect 7196 14000 7248 14006
rect 7196 13942 7248 13948
rect 7288 14000 7340 14006
rect 7288 13942 7340 13948
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 5644 12238 5672 12718
rect 5828 12374 5856 13806
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6472 12374 6500 12718
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 5816 12368 5868 12374
rect 5816 12310 5868 12316
rect 6460 12368 6512 12374
rect 6460 12310 6512 12316
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 3514 12064 3570 12073
rect 3514 11999 3570 12008
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2792 10606 2820 11154
rect 3068 11150 3096 11698
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3160 10810 3188 11630
rect 5092 11354 5120 11630
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3988 10606 4016 11154
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3988 10062 4016 10542
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 2778 9888 2834 9897
rect 2778 9823 2834 9832
rect 388 9172 440 9178
rect 388 9114 440 9120
rect 400 800 428 9114
rect 2792 8634 2820 9823
rect 3988 9586 4016 9998
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 9042 3004 9318
rect 3252 9110 3280 9454
rect 3240 9104 3292 9110
rect 3240 9046 3292 9052
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2884 8922 2912 8978
rect 3056 8968 3108 8974
rect 2884 8894 3004 8922
rect 3056 8910 3108 8916
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1872 6905 1900 8366
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 1858 6896 1914 6905
rect 1858 6831 1914 6840
rect 2688 6248 2740 6254
rect 2686 6216 2688 6225
rect 2740 6216 2742 6225
rect 2686 6151 2742 6160
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2792 5545 2820 6054
rect 2884 5574 2912 7890
rect 2872 5568 2924 5574
rect 2778 5536 2834 5545
rect 2872 5510 2924 5516
rect 2778 5471 2834 5480
rect 2976 5370 3004 8894
rect 3068 7886 3096 8910
rect 3988 8498 4016 9522
rect 4080 8634 4108 10406
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3160 7818 3188 8366
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 3054 7712 3110 7721
rect 3054 7647 3110 7656
rect 3068 7002 3096 7647
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 3160 6322 3188 7278
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2872 5160 2924 5166
rect 2700 5120 2872 5148
rect 2700 4690 2728 5120
rect 2872 5102 2924 5108
rect 3252 4758 3280 7890
rect 3988 7410 4016 8434
rect 4080 8022 4108 8570
rect 4356 8022 4384 9998
rect 4068 8016 4120 8022
rect 4068 7958 4120 7964
rect 4344 8016 4396 8022
rect 4344 7958 4396 7964
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3988 6866 4016 7346
rect 4252 7268 4304 7274
rect 4252 7210 4304 7216
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4172 5166 4200 6802
rect 4264 5778 4292 7210
rect 4448 7206 4476 11018
rect 4724 9110 4752 11086
rect 5460 10674 5488 11630
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4356 5846 4384 6734
rect 4448 6254 4476 7142
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4160 5160 4212 5166
rect 4212 5108 4384 5114
rect 4160 5102 4384 5108
rect 4172 5086 4384 5102
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 2700 4078 2728 4626
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 3976 4072 4028 4078
rect 4080 4049 4108 4626
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 3976 4014 4028 4020
rect 4066 4040 4122 4049
rect 1214 3768 1270 3777
rect 3988 3738 4016 4014
rect 4066 3975 4122 3984
rect 1214 3703 1270 3712
rect 3976 3732 4028 3738
rect 1228 800 1256 3703
rect 3976 3674 4028 3680
rect 3790 3496 3846 3505
rect 3790 3431 3846 3440
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 2056 800 2084 2450
rect 2976 800 3004 2450
rect 3424 1352 3476 1358
rect 3424 1294 3476 1300
rect 3436 1193 3464 1294
rect 3422 1184 3478 1193
rect 3422 1119 3478 1128
rect 3804 800 3832 3431
rect 4066 3360 4122 3369
rect 4172 3346 4200 4422
rect 4122 3318 4200 3346
rect 4066 3295 4122 3304
rect 4356 2446 4384 5086
rect 4540 4146 4568 8978
rect 5092 7954 5120 10202
rect 5552 9042 5580 11018
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5644 8634 5672 8978
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5368 6254 5396 8366
rect 5644 7954 5672 8570
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 4816 5778 4844 6190
rect 5552 5846 5580 6598
rect 5644 6322 5672 7482
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5736 5778 5764 6802
rect 6380 6322 6408 12242
rect 6564 10062 6592 12582
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6840 11150 6868 12174
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6932 11286 6960 11630
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6656 10130 6684 10746
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6564 6882 6592 9998
rect 6748 9654 6776 10542
rect 7024 10198 7052 12650
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 7116 10810 7144 12106
rect 7208 11898 7236 13942
rect 7392 13938 7420 14350
rect 7576 13938 7604 14894
rect 8128 14550 8156 15574
rect 8588 15570 8616 18835
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8588 15162 8616 15506
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8312 12850 8340 13806
rect 10152 13394 10180 15846
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10336 13802 10364 15438
rect 10428 14822 10456 15506
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 10428 13462 10456 14758
rect 10520 14482 10548 18835
rect 11137 17436 11433 17456
rect 11193 17434 11217 17436
rect 11273 17434 11297 17436
rect 11353 17434 11377 17436
rect 11215 17382 11217 17434
rect 11279 17382 11291 17434
rect 11353 17382 11355 17434
rect 11193 17380 11217 17382
rect 11273 17380 11297 17382
rect 11353 17380 11377 17382
rect 11137 17360 11433 17380
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11716 16658 11744 17138
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11137 16348 11433 16368
rect 11193 16346 11217 16348
rect 11273 16346 11297 16348
rect 11353 16346 11377 16348
rect 11215 16294 11217 16346
rect 11279 16294 11291 16346
rect 11353 16294 11355 16346
rect 11193 16292 11217 16294
rect 11273 16292 11297 16294
rect 11353 16292 11377 16294
rect 11137 16272 11433 16292
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10968 14884 11020 14890
rect 10968 14826 11020 14832
rect 10980 14618 11008 14826
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 11072 14074 11100 15302
rect 11137 15260 11433 15280
rect 11193 15258 11217 15260
rect 11273 15258 11297 15260
rect 11353 15258 11377 15260
rect 11215 15206 11217 15258
rect 11279 15206 11291 15258
rect 11353 15206 11355 15258
rect 11193 15204 11217 15206
rect 11273 15204 11297 15206
rect 11353 15204 11377 15206
rect 11137 15184 11433 15204
rect 11716 14958 11744 16594
rect 12164 16040 12216 16046
rect 12164 15982 12216 15988
rect 12176 15570 12204 15982
rect 12348 15972 12400 15978
rect 12348 15914 12400 15920
rect 12360 15706 12388 15914
rect 12348 15700 12400 15706
rect 12348 15642 12400 15648
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 12452 15094 12480 18835
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12544 15366 12572 16594
rect 13096 16250 13124 17070
rect 14292 16726 14320 18835
rect 16224 17338 16252 18835
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 14280 16720 14332 16726
rect 14280 16662 14332 16668
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 12716 16040 12768 16046
rect 12636 16000 12716 16028
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11716 14414 11744 14894
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11137 14172 11433 14192
rect 11193 14170 11217 14172
rect 11273 14170 11297 14172
rect 11353 14170 11377 14172
rect 11215 14118 11217 14170
rect 11279 14118 11291 14170
rect 11353 14118 11355 14170
rect 11193 14116 11217 14118
rect 11273 14116 11297 14118
rect 11353 14116 11377 14118
rect 11137 14096 11433 14116
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12360 13938 12388 14010
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 10966 13560 11022 13569
rect 10966 13495 11022 13504
rect 10416 13456 10468 13462
rect 10416 13398 10468 13404
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 7300 12102 7328 12786
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7484 12306 7512 12718
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7300 10470 7328 12038
rect 7484 11082 7512 12242
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7576 11762 7604 12106
rect 7944 11762 7972 12174
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7576 10810 7604 11698
rect 8220 11694 8248 12038
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 7668 9518 7696 10406
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6656 7342 6684 7754
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6472 6866 6592 6882
rect 6656 6866 6684 7278
rect 6460 6860 6592 6866
rect 6512 6854 6592 6860
rect 6644 6860 6696 6866
rect 6460 6802 6512 6808
rect 6644 6802 6696 6808
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 6380 5370 6408 6258
rect 6920 6248 6972 6254
rect 6840 6208 6920 6236
rect 6736 5840 6788 5846
rect 6840 5794 6868 6208
rect 6920 6190 6972 6196
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6788 5788 6868 5794
rect 6736 5782 6868 5788
rect 6748 5766 6868 5782
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5368 4758 5396 5102
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 5736 4078 5764 5034
rect 6380 4826 6408 5306
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 5814 4720 5870 4729
rect 5814 4655 5816 4664
rect 5868 4655 5870 4664
rect 5816 4626 5868 4632
rect 6840 4214 6868 5766
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 6932 4690 6960 5578
rect 7024 5370 7052 6054
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 7116 4622 7144 6054
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 6828 4208 6880 4214
rect 6656 4156 6828 4162
rect 6656 4150 6880 4156
rect 6656 4134 6868 4150
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 4710 3088 4766 3097
rect 5000 3058 5028 3470
rect 5368 3466 5396 4014
rect 6656 3670 6684 4134
rect 6932 4026 6960 4218
rect 7208 4146 7236 9454
rect 7484 9042 7512 9454
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7300 5778 7328 6054
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7300 5166 7328 5714
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 6840 3998 6960 4026
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 3670 6776 3878
rect 6644 3664 6696 3670
rect 6366 3632 6422 3641
rect 6644 3606 6696 3612
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6366 3567 6422 3576
rect 6460 3596 6512 3602
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 4710 3023 4766 3032
rect 4988 3052 5040 3058
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4724 800 4752 3023
rect 4988 2994 5040 3000
rect 5552 2514 5580 3334
rect 5630 2952 5686 2961
rect 5630 2887 5686 2896
rect 5908 2916 5960 2922
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5644 1034 5672 2887
rect 5908 2858 5960 2864
rect 5920 2514 5948 2858
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 5552 1006 5672 1034
rect 5552 800 5580 1006
rect 6380 800 6408 3567
rect 6460 3538 6512 3544
rect 6472 3194 6500 3538
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6564 3126 6592 3470
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6840 2990 6868 3998
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6932 3058 6960 3878
rect 7392 3602 7420 4558
rect 7760 4146 7788 6734
rect 8036 5778 8064 11630
rect 8760 10600 8812 10606
rect 8758 10568 8760 10577
rect 8812 10568 8814 10577
rect 8758 10503 8814 10512
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8208 8968 8260 8974
rect 8260 8916 8340 8922
rect 8208 8910 8340 8916
rect 8220 8894 8340 8910
rect 8312 7954 8340 8894
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 8498 8432 8774
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8680 8430 8708 9318
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8680 7410 8708 8366
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8772 7410 8800 7822
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 7838 5264 7894 5273
rect 7838 5199 7894 5208
rect 7852 5166 7880 5199
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7944 5030 7972 5714
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7484 3466 7512 4014
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 7472 3460 7524 3466
rect 7472 3402 7524 3408
rect 7576 3194 7604 3946
rect 7944 3602 7972 4966
rect 8036 4282 8064 5714
rect 8128 4690 8156 7346
rect 8772 6934 8800 7346
rect 8760 6928 8812 6934
rect 8760 6870 8812 6876
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8220 5166 8248 5850
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8404 5234 8432 5646
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8116 4684 8168 4690
rect 8116 4626 8168 4632
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 8024 3460 8076 3466
rect 8024 3402 8076 3408
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7852 3058 7880 3402
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8036 2990 8064 3402
rect 8128 3074 8156 4626
rect 8220 3534 8248 5102
rect 8404 4758 8432 5170
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 8588 3602 8616 6802
rect 8956 5914 8984 12854
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9048 11218 9076 11630
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 9232 10577 9260 12718
rect 9324 12374 9352 12718
rect 9312 12368 9364 12374
rect 9312 12310 9364 12316
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9692 10810 9720 10950
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9218 10568 9274 10577
rect 9218 10503 9274 10512
rect 9680 10056 9732 10062
rect 9600 10004 9680 10010
rect 9600 9998 9732 10004
rect 9600 9982 9720 9998
rect 9600 9330 9628 9982
rect 9680 9376 9732 9382
rect 9600 9324 9680 9330
rect 9600 9318 9732 9324
rect 9600 9302 9720 9318
rect 9600 9110 9628 9302
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9784 7478 9812 13330
rect 10152 13190 10180 13330
rect 10782 13288 10838 13297
rect 10782 13223 10838 13232
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9876 12345 9904 12378
rect 9862 12336 9918 12345
rect 10796 12306 10824 13223
rect 9862 12271 9918 12280
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10980 12238 11008 13495
rect 11072 13326 11100 13806
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11072 12782 11100 13262
rect 11137 13084 11433 13104
rect 11193 13082 11217 13084
rect 11273 13082 11297 13084
rect 11353 13082 11377 13084
rect 11215 13030 11217 13082
rect 11279 13030 11291 13082
rect 11353 13030 11355 13082
rect 11193 13028 11217 13030
rect 11273 13028 11297 13030
rect 11353 13028 11377 13030
rect 11137 13008 11433 13028
rect 11532 12782 11560 13806
rect 12544 13802 12572 14826
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 11060 12776 11112 12782
rect 11520 12776 11572 12782
rect 11060 12718 11112 12724
rect 11440 12736 11520 12764
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 11164 12084 11192 12378
rect 11256 12220 11284 12650
rect 11440 12374 11468 12736
rect 11520 12718 11572 12724
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11428 12232 11480 12238
rect 11256 12192 11428 12220
rect 11428 12174 11480 12180
rect 11072 12056 11192 12084
rect 11072 11694 11100 12056
rect 11137 11996 11433 12016
rect 11193 11994 11217 11996
rect 11273 11994 11297 11996
rect 11353 11994 11377 11996
rect 11215 11942 11217 11994
rect 11279 11942 11291 11994
rect 11353 11942 11355 11994
rect 11193 11940 11217 11942
rect 11273 11940 11297 11942
rect 11353 11940 11377 11942
rect 11137 11920 11433 11940
rect 11532 11762 11560 12242
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11060 11688 11112 11694
rect 11256 11665 11284 11698
rect 11336 11688 11388 11694
rect 11060 11630 11112 11636
rect 11242 11656 11298 11665
rect 10782 11248 10838 11257
rect 10782 11183 10784 11192
rect 10836 11183 10838 11192
rect 10968 11212 11020 11218
rect 10784 11154 10836 11160
rect 11072 11200 11100 11630
rect 11336 11630 11388 11636
rect 11242 11591 11298 11600
rect 11348 11286 11376 11630
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11020 11172 11100 11200
rect 10968 11154 11020 11160
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9876 9722 9904 10542
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10060 10130 10088 10406
rect 10796 10266 10824 11154
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10048 10124 10100 10130
rect 10048 10066 10100 10072
rect 10888 10062 10916 10950
rect 11137 10908 11433 10928
rect 11193 10906 11217 10908
rect 11273 10906 11297 10908
rect 11353 10906 11377 10908
rect 11215 10854 11217 10906
rect 11279 10854 11291 10906
rect 11353 10854 11355 10906
rect 11193 10852 11217 10854
rect 11273 10852 11297 10854
rect 11353 10852 11377 10854
rect 11137 10832 11433 10852
rect 11610 10840 11666 10849
rect 11610 10775 11666 10784
rect 11624 10606 11652 10775
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 10980 10470 11008 10542
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9692 6458 9720 7278
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8956 5166 8984 5850
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8680 4010 8708 4422
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 8668 4004 8720 4010
rect 8668 3946 8720 3952
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8128 3058 8248 3074
rect 8128 3052 8260 3058
rect 8128 3046 8208 3052
rect 8208 2994 8260 3000
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 6840 2582 6868 2926
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 6828 2576 6880 2582
rect 6828 2518 6880 2524
rect 7300 800 7328 2790
rect 8128 800 8156 2926
rect 8680 2582 8708 3946
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 9048 800 9076 4082
rect 9140 3942 9168 5102
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9140 3398 9168 3878
rect 9784 3777 9812 7414
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9968 6866 9996 7210
rect 10060 6934 10088 8366
rect 10244 7886 10272 9862
rect 10980 9586 11008 10406
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11137 9820 11433 9840
rect 11193 9818 11217 9820
rect 11273 9818 11297 9820
rect 11353 9818 11377 9820
rect 11215 9766 11217 9818
rect 11279 9766 11291 9818
rect 11353 9766 11355 9818
rect 11193 9764 11217 9766
rect 11273 9764 11297 9766
rect 11353 9764 11377 9766
rect 11137 9744 11433 9764
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11532 9518 11560 9862
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 10336 6798 10364 7890
rect 10612 6866 10640 8978
rect 11072 8974 11100 9454
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10796 8090 10824 8910
rect 11137 8732 11433 8752
rect 11193 8730 11217 8732
rect 11273 8730 11297 8732
rect 11353 8730 11377 8732
rect 11215 8678 11217 8730
rect 11279 8678 11291 8730
rect 11353 8678 11355 8730
rect 11193 8676 11217 8678
rect 11273 8676 11297 8678
rect 11353 8676 11377 8678
rect 11137 8656 11433 8676
rect 11532 8634 11560 9454
rect 11624 9058 11652 10066
rect 11716 9994 11744 13738
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11992 12782 12020 13262
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11808 9382 11836 10202
rect 11900 10130 11928 12242
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12176 10674 12204 11086
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12072 10532 12124 10538
rect 12072 10474 12124 10480
rect 12084 10130 12112 10474
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11796 9104 11848 9110
rect 11624 9052 11796 9058
rect 11624 9046 11848 9052
rect 11624 9030 11836 9046
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11624 8430 11652 9030
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 10152 6322 10180 6666
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10244 6254 10272 6598
rect 10612 6254 10640 6802
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10704 4185 10732 7890
rect 10888 5166 10916 8366
rect 11164 8022 11192 8366
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11137 7644 11433 7664
rect 11193 7642 11217 7644
rect 11273 7642 11297 7644
rect 11353 7642 11377 7644
rect 11215 7590 11217 7642
rect 11279 7590 11291 7642
rect 11353 7590 11355 7642
rect 11193 7588 11217 7590
rect 11273 7588 11297 7590
rect 11353 7588 11377 7590
rect 11137 7568 11433 7588
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10980 5642 11008 7278
rect 11137 6556 11433 6576
rect 11193 6554 11217 6556
rect 11273 6554 11297 6556
rect 11353 6554 11377 6556
rect 11215 6502 11217 6554
rect 11279 6502 11291 6554
rect 11353 6502 11355 6554
rect 11193 6500 11217 6502
rect 11273 6500 11297 6502
rect 11353 6500 11377 6502
rect 11137 6480 11433 6500
rect 11808 5778 11836 7686
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 11900 6866 11928 7210
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11992 6322 12020 6734
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 12084 6118 12112 9930
rect 12176 9586 12204 10610
rect 12268 10266 12296 13330
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12360 12374 12388 13262
rect 12636 12986 12664 16000
rect 12716 15982 12768 15988
rect 13832 15570 13860 16662
rect 14384 16046 14412 17274
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 15304 16726 15332 17002
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 15292 16720 15344 16726
rect 15292 16662 15344 16668
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12728 14074 12756 14894
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13004 14074 13032 14350
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 12348 11824 12400 11830
rect 12346 11792 12348 11801
rect 12400 11792 12402 11801
rect 12346 11727 12402 11736
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12452 11014 12480 11698
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12346 9072 12402 9081
rect 12346 9007 12348 9016
rect 12400 9007 12402 9016
rect 12348 8978 12400 8984
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10876 5160 10928 5166
rect 10980 5137 11008 5578
rect 11137 5468 11433 5488
rect 11193 5466 11217 5468
rect 11273 5466 11297 5468
rect 11353 5466 11377 5468
rect 11215 5414 11217 5466
rect 11279 5414 11291 5466
rect 11353 5414 11355 5466
rect 11193 5412 11217 5414
rect 11273 5412 11297 5414
rect 11353 5412 11377 5414
rect 11137 5392 11433 5412
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10876 5102 10928 5108
rect 10966 5128 11022 5137
rect 10966 5063 11022 5072
rect 11072 4214 11100 5170
rect 12176 4690 12204 6802
rect 12268 5234 12296 8910
rect 12544 6322 12572 12582
rect 12728 11830 12756 13806
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12912 13138 12940 13194
rect 13084 13184 13136 13190
rect 12912 13110 13032 13138
rect 13084 13126 13136 13132
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12912 11937 12940 12174
rect 13004 12102 13032 13110
rect 13096 12782 13124 13126
rect 13280 12850 13308 13262
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 12898 11928 12954 11937
rect 12898 11863 12954 11872
rect 12716 11824 12768 11830
rect 13096 11778 13124 12106
rect 13372 12102 13400 12718
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 12716 11766 12768 11772
rect 13004 11750 13124 11778
rect 13004 11642 13032 11750
rect 12820 11614 13032 11642
rect 12820 11558 12848 11614
rect 12808 11552 12860 11558
rect 13188 11529 13216 11834
rect 13280 11801 13308 11834
rect 13266 11792 13322 11801
rect 13266 11727 13322 11736
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13268 11688 13320 11694
rect 13372 11665 13400 11698
rect 13268 11630 13320 11636
rect 13358 11656 13414 11665
rect 12808 11494 12860 11500
rect 13174 11520 13230 11529
rect 13174 11455 13230 11464
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13188 10470 13216 11290
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 12716 9512 12768 9518
rect 12716 9454 12768 9460
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 12728 8022 12756 9454
rect 12716 8016 12768 8022
rect 12622 7984 12678 7993
rect 12716 7958 12768 7964
rect 12622 7919 12624 7928
rect 12676 7919 12678 7928
rect 12624 7890 12676 7896
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12636 6202 12664 7890
rect 13004 7410 13032 9454
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13096 6662 13124 6734
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12532 6180 12584 6186
rect 12636 6174 12848 6202
rect 12532 6122 12584 6128
rect 12544 6066 12572 6122
rect 12452 6038 12572 6066
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12452 5778 12480 6038
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12176 4593 12204 4626
rect 12162 4584 12218 4593
rect 12162 4519 12218 4528
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11137 4380 11433 4400
rect 11193 4378 11217 4380
rect 11273 4378 11297 4380
rect 11353 4378 11377 4380
rect 11215 4326 11217 4378
rect 11279 4326 11291 4378
rect 11353 4326 11355 4378
rect 11193 4324 11217 4326
rect 11273 4324 11297 4326
rect 11353 4324 11377 4326
rect 11137 4304 11433 4324
rect 11992 4282 12020 4422
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11060 4208 11112 4214
rect 9954 4176 10010 4185
rect 9954 4111 10010 4120
rect 10690 4176 10746 4185
rect 11060 4150 11112 4156
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 10690 4111 10746 4120
rect 9968 4010 9996 4111
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9770 3768 9826 3777
rect 9770 3703 9826 3712
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9876 800 9904 2994
rect 10796 800 10824 3470
rect 11137 3292 11433 3312
rect 11193 3290 11217 3292
rect 11273 3290 11297 3292
rect 11353 3290 11377 3292
rect 11215 3238 11217 3290
rect 11279 3238 11291 3290
rect 11353 3238 11355 3290
rect 11193 3236 11217 3238
rect 11273 3236 11297 3238
rect 11353 3236 11377 3238
rect 11137 3216 11433 3236
rect 11137 2204 11433 2224
rect 11193 2202 11217 2204
rect 11273 2202 11297 2204
rect 11353 2202 11377 2204
rect 11215 2150 11217 2202
rect 11279 2150 11291 2202
rect 11353 2150 11355 2202
rect 11193 2148 11217 2150
rect 11273 2148 11297 2150
rect 11353 2148 11377 2150
rect 11137 2128 11433 2148
rect 11624 800 11652 4150
rect 12360 2514 12388 5714
rect 12452 5574 12480 5714
rect 12636 5710 12664 6054
rect 12728 5914 12756 6054
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12452 4758 12480 5510
rect 12544 5370 12572 5646
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12440 4752 12492 4758
rect 12820 4729 12848 6174
rect 13096 5166 13124 6598
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12440 4694 12492 4700
rect 12806 4720 12862 4729
rect 13188 4690 13216 9998
rect 12806 4655 12862 4664
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12452 3534 12480 4490
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12348 2508 12400 2514
rect 12348 2450 12400 2456
rect 12452 800 12480 3470
rect 12728 1970 12756 3606
rect 12820 3602 12848 4558
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12820 2446 12848 3538
rect 13004 3194 13032 3606
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13096 3194 13124 3538
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13188 3126 13216 4014
rect 13280 4010 13308 11630
rect 13358 11591 13414 11600
rect 13372 10130 13400 11591
rect 13464 11082 13492 13262
rect 13636 13252 13688 13258
rect 13636 13194 13688 13200
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13556 10010 13584 12038
rect 13648 11762 13676 13194
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13740 10198 13768 13806
rect 14200 13802 14228 14214
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14016 12102 14044 12718
rect 14660 12646 14688 13330
rect 15212 12714 15240 15982
rect 15304 15978 15332 16662
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15304 15434 15332 15914
rect 15488 15570 15516 16050
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15488 14482 15516 15506
rect 16316 15162 16344 16118
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 16500 14958 16528 16526
rect 16592 15978 16620 16934
rect 16684 16658 16712 17138
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17684 17060 17736 17066
rect 17684 17002 17736 17008
rect 17696 16726 17724 17002
rect 17684 16720 17736 16726
rect 17684 16662 17736 16668
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 16684 15570 16712 16594
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15384 13796 15436 13802
rect 15384 13738 15436 13744
rect 15396 13462 15424 13738
rect 16592 13569 16620 14894
rect 16684 14482 16712 15506
rect 16960 15162 16988 16594
rect 17224 15972 17276 15978
rect 17224 15914 17276 15920
rect 17236 15570 17264 15914
rect 17972 15638 18000 17070
rect 18156 16794 18184 18835
rect 20088 17338 20116 18835
rect 20076 17332 20128 17338
rect 20076 17274 20128 17280
rect 18420 17128 18472 17134
rect 18420 17070 18472 17076
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18432 16590 18460 17070
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18236 16448 18288 16454
rect 18236 16390 18288 16396
rect 18248 16046 18276 16390
rect 18236 16040 18288 16046
rect 18236 15982 18288 15988
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 17960 14544 18012 14550
rect 17960 14486 18012 14492
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16578 13560 16634 13569
rect 16578 13495 16634 13504
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15304 13297 15332 13330
rect 15290 13288 15346 13297
rect 15290 13223 15346 13232
rect 16684 12866 16712 14418
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17144 13462 17172 14350
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 17972 13394 18000 14486
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 16592 12838 16712 12866
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 14016 11218 14044 12038
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14384 11286 14412 11766
rect 15028 11762 15056 12242
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 14464 11620 14516 11626
rect 14464 11562 14516 11568
rect 14556 11620 14608 11626
rect 14556 11562 14608 11568
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13820 10056 13872 10062
rect 13452 9988 13504 9994
rect 13556 9982 13768 10010
rect 13820 9998 13872 10004
rect 13452 9930 13504 9936
rect 13464 9722 13492 9930
rect 13740 9926 13768 9982
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13740 9518 13768 9862
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13832 9450 13860 9998
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 13372 7342 13400 8366
rect 13556 7954 13584 8502
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13740 7546 13768 8978
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13832 7886 13860 8774
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13464 7206 13492 7278
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13464 5273 13492 7142
rect 14108 6866 14136 11154
rect 14476 10674 14504 11562
rect 14568 11257 14596 11562
rect 14936 11286 14964 11630
rect 14924 11280 14976 11286
rect 14554 11248 14610 11257
rect 14924 11222 14976 11228
rect 14554 11183 14610 11192
rect 15028 10742 15056 11698
rect 15120 11234 15148 12038
rect 15396 11762 15424 12038
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15120 11206 15240 11234
rect 15212 11150 15240 11206
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 15120 10198 15148 11086
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15108 10192 15160 10198
rect 15108 10134 15160 10140
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 14280 9104 14332 9110
rect 14280 9046 14332 9052
rect 14292 8634 14320 9046
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14292 7750 14320 8570
rect 14660 8430 14688 9386
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14660 7342 14688 7890
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 13832 5914 13860 6802
rect 14476 6730 14504 7278
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13450 5264 13506 5273
rect 13740 5234 13768 5510
rect 13450 5199 13506 5208
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13556 4146 13584 5102
rect 13740 5030 13768 5170
rect 14108 5098 14136 6598
rect 14096 5092 14148 5098
rect 14096 5034 14148 5040
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13636 4752 13688 4758
rect 13636 4694 13688 4700
rect 13648 4282 13676 4694
rect 13740 4690 13768 4966
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14016 4282 14044 4558
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 13268 4004 13320 4010
rect 13268 3946 13320 3952
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13280 3398 13308 3946
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 13464 3058 13492 3946
rect 14200 3738 14228 4014
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13740 2990 13768 3470
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 13924 2990 13952 3334
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 12912 2514 12940 2858
rect 12900 2508 12952 2514
rect 12900 2450 12952 2456
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 12716 1964 12768 1970
rect 12716 1906 12768 1912
rect 13360 1964 13412 1970
rect 13360 1906 13412 1912
rect 13372 800 13400 1906
rect 14200 800 14228 3674
rect 14476 2038 14504 6666
rect 14936 5370 14964 7482
rect 15028 7410 15056 10066
rect 15304 9654 15332 10542
rect 15396 10198 15424 11698
rect 15764 11558 15792 12718
rect 16592 12646 16620 12838
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15384 10192 15436 10198
rect 15384 10134 15436 10140
rect 15292 9648 15344 9654
rect 15292 9590 15344 9596
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15396 7750 15424 9454
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15108 6860 15160 6866
rect 15108 6802 15160 6808
rect 15016 6180 15068 6186
rect 15016 6122 15068 6128
rect 15028 5846 15056 6122
rect 15016 5840 15068 5846
rect 15016 5782 15068 5788
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 14738 3360 14794 3369
rect 14738 3295 14794 3304
rect 14752 2990 14780 3295
rect 14740 2984 14792 2990
rect 14740 2926 14792 2932
rect 14464 2032 14516 2038
rect 14464 1974 14516 1980
rect 15120 800 15148 6802
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15212 5166 15240 5714
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15304 5234 15332 5578
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15212 4826 15240 5102
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15396 4622 15424 5646
rect 15488 5574 15516 6190
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15580 5030 15608 8434
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15672 7206 15700 7686
rect 15764 7206 15792 10406
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15856 9586 15884 10066
rect 16040 10010 16068 11154
rect 16132 11082 16160 12310
rect 16684 12306 16712 12718
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16408 12170 16620 12186
rect 16396 12164 16620 12170
rect 16448 12158 16620 12164
rect 16396 12106 16448 12112
rect 16394 11928 16450 11937
rect 16394 11863 16450 11872
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 16132 10130 16160 11018
rect 16224 10452 16252 11630
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16316 10606 16344 11494
rect 16408 10742 16436 11863
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16396 10464 16448 10470
rect 16224 10424 16396 10452
rect 16396 10406 16448 10412
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 16040 9982 16160 10010
rect 16028 9920 16080 9926
rect 16028 9862 16080 9868
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15948 8090 15976 8774
rect 16040 8430 16068 9862
rect 16132 8838 16160 9982
rect 16408 9042 16436 10406
rect 16592 9518 16620 12158
rect 16672 10736 16724 10742
rect 16672 10678 16724 10684
rect 16684 9586 16712 10678
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 17052 9110 17080 13330
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17236 12986 17264 13194
rect 18156 12986 18184 13874
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17604 12782 17632 12854
rect 17592 12776 17644 12782
rect 17592 12718 17644 12724
rect 17604 12306 17632 12718
rect 17774 12336 17830 12345
rect 17592 12300 17644 12306
rect 17774 12271 17776 12280
rect 17592 12242 17644 12248
rect 17828 12271 17830 12280
rect 17776 12242 17828 12248
rect 17500 11620 17552 11626
rect 17500 11562 17552 11568
rect 17512 11014 17540 11562
rect 18248 11286 18276 13806
rect 18340 13802 18368 15982
rect 18432 14958 18460 16526
rect 18616 16250 18644 17070
rect 20088 16658 20116 17274
rect 21318 16892 21614 16912
rect 21374 16890 21398 16892
rect 21454 16890 21478 16892
rect 21534 16890 21558 16892
rect 21396 16838 21398 16890
rect 21460 16838 21472 16890
rect 21534 16838 21536 16890
rect 21374 16836 21398 16838
rect 21454 16836 21478 16838
rect 21534 16836 21558 16838
rect 21318 16816 21614 16836
rect 20076 16652 20128 16658
rect 20076 16594 20128 16600
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 20628 16040 20680 16046
rect 20680 16000 20760 16028
rect 20628 15982 20680 15988
rect 19524 15972 19576 15978
rect 19524 15914 19576 15920
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18432 13938 18460 14894
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18328 13796 18380 13802
rect 18328 13738 18380 13744
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17512 9654 17540 10950
rect 18432 10810 18460 13874
rect 18800 13462 18828 14894
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19444 14482 19472 14758
rect 19536 14482 19564 15914
rect 19708 15564 19760 15570
rect 19708 15506 19760 15512
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19536 14090 19564 14418
rect 19444 14062 19564 14090
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18892 12714 18920 13466
rect 19076 13297 19104 13466
rect 19444 13433 19472 14062
rect 19430 13424 19486 13433
rect 19430 13359 19486 13368
rect 19524 13388 19576 13394
rect 19062 13288 19118 13297
rect 19062 13223 19118 13232
rect 19444 12714 19472 13359
rect 19524 13330 19576 13336
rect 18788 12708 18840 12714
rect 18788 12650 18840 12656
rect 18880 12708 18932 12714
rect 18880 12650 18932 12656
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 18800 11626 18828 12650
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18892 11937 18920 12378
rect 19352 12374 19380 12582
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 18878 11928 18934 11937
rect 18878 11863 18934 11872
rect 18788 11620 18840 11626
rect 18788 11562 18840 11568
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 18786 11520 18842 11529
rect 18786 11455 18842 11464
rect 18800 11286 18828 11455
rect 18788 11280 18840 11286
rect 18788 11222 18840 11228
rect 19352 11218 19380 11562
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19248 11144 19300 11150
rect 19300 11092 19380 11098
rect 19248 11086 19380 11092
rect 19260 11070 19380 11086
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 19352 10606 19380 11070
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19248 10532 19300 10538
rect 19248 10474 19300 10480
rect 18972 10464 19024 10470
rect 19064 10464 19116 10470
rect 19024 10424 19064 10452
rect 18972 10406 19024 10412
rect 19064 10406 19116 10412
rect 19260 10266 19288 10474
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19444 10130 19472 10406
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17500 9648 17552 9654
rect 17500 9590 17552 9596
rect 17604 9466 17632 9998
rect 18432 9518 18460 10066
rect 19340 10056 19392 10062
rect 19338 10024 19340 10033
rect 19392 10024 19394 10033
rect 19338 9959 19394 9968
rect 17512 9438 17632 9466
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15764 6798 15792 7142
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15764 5778 15792 6734
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15672 5658 15700 5714
rect 15672 5630 15792 5658
rect 15764 5166 15792 5630
rect 15856 5352 15884 7822
rect 15948 7342 15976 8026
rect 16132 7954 16160 8774
rect 16500 8090 16528 8910
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 16500 7410 16528 8026
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 16396 7200 16448 7206
rect 16132 7160 16396 7188
rect 16132 6934 16160 7160
rect 16396 7142 16448 7148
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16316 6322 16344 6734
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 15856 5324 15976 5352
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 15672 4842 15700 4966
rect 15580 4814 15700 4842
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15580 4486 15608 4814
rect 15764 4554 15792 5102
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15580 4298 15608 4422
rect 15212 4270 15608 4298
rect 15212 4146 15240 4270
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15304 3913 15332 4014
rect 15290 3904 15346 3913
rect 15290 3839 15346 3848
rect 15580 3534 15608 4270
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15948 800 15976 5324
rect 16224 4826 16252 6258
rect 16592 6254 16620 7822
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 16764 7336 16816 7342
rect 16684 7296 16764 7324
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16684 6118 16712 7296
rect 16764 7278 16816 7284
rect 17144 6390 17172 7346
rect 17132 6384 17184 6390
rect 17132 6326 17184 6332
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16316 4690 16344 5646
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16028 4548 16080 4554
rect 16028 4490 16080 4496
rect 16040 4010 16068 4490
rect 16028 4004 16080 4010
rect 16028 3946 16080 3952
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16040 3466 16068 3674
rect 16316 3602 16344 4626
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16316 2854 16344 3402
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 16408 2446 16436 5714
rect 17512 5574 17540 9438
rect 18340 9382 18368 9454
rect 18328 9376 18380 9382
rect 18328 9318 18380 9324
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 18696 9104 18748 9110
rect 17958 9072 18014 9081
rect 18696 9046 18748 9052
rect 17958 9007 18014 9016
rect 18512 9036 18564 9042
rect 17776 8968 17828 8974
rect 17774 8936 17776 8945
rect 17828 8936 17830 8945
rect 17972 8906 18000 9007
rect 18512 8978 18564 8984
rect 17774 8871 17830 8880
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 18524 8430 18552 8978
rect 18708 8430 18736 9046
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 17604 7954 17632 8298
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16684 5166 16712 5306
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16684 4078 16712 4558
rect 16868 4078 16896 4558
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 16592 2689 16620 2790
rect 16578 2680 16634 2689
rect 16578 2615 16634 2624
rect 16684 2446 16712 4014
rect 16868 3602 16896 4014
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16960 2990 16988 4762
rect 17236 4078 17264 5102
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17236 3602 17264 4014
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17236 3369 17264 3538
rect 17512 3534 17540 5510
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17222 3360 17278 3369
rect 17222 3295 17278 3304
rect 17592 3120 17644 3126
rect 17592 3062 17644 3068
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 16776 2825 16804 2926
rect 17316 2916 17368 2922
rect 17316 2858 17368 2864
rect 16762 2816 16818 2825
rect 16762 2751 16818 2760
rect 17328 2514 17356 2858
rect 17604 2514 17632 3062
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 16396 2440 16448 2446
rect 16396 2382 16448 2388
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 16408 2106 16436 2382
rect 16396 2100 16448 2106
rect 16396 2042 16448 2048
rect 16856 2032 16908 2038
rect 16856 1974 16908 1980
rect 16868 800 16896 1974
rect 17696 800 17724 8026
rect 17868 8016 17920 8022
rect 17866 7984 17868 7993
rect 17920 7984 17922 7993
rect 17866 7919 17922 7928
rect 18708 7886 18736 8366
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17972 6730 18000 7210
rect 18064 6934 18092 7822
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18800 6934 18828 7278
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 18788 6928 18840 6934
rect 18788 6870 18840 6876
rect 19260 6798 19288 7822
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 19352 6662 19380 9318
rect 19444 8956 19472 10066
rect 19536 9586 19564 13330
rect 19628 12918 19656 15302
rect 19616 12912 19668 12918
rect 19616 12854 19668 12860
rect 19720 12374 19748 15506
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19812 13394 19840 14758
rect 20732 14550 20760 16000
rect 21180 15972 21232 15978
rect 21180 15914 21232 15920
rect 21192 14958 21220 15914
rect 21318 15804 21614 15824
rect 21374 15802 21398 15804
rect 21454 15802 21478 15804
rect 21534 15802 21558 15804
rect 21396 15750 21398 15802
rect 21460 15750 21472 15802
rect 21534 15750 21536 15802
rect 21374 15748 21398 15750
rect 21454 15748 21478 15750
rect 21534 15748 21558 15750
rect 21318 15728 21614 15748
rect 22020 15638 22048 18835
rect 22560 17060 22612 17066
rect 22560 17002 22612 17008
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22204 15978 22232 16934
rect 22572 16726 22600 17002
rect 23952 16794 23980 18835
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 24032 17128 24084 17134
rect 24032 17070 24084 17076
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 23940 16788 23992 16794
rect 23940 16730 23992 16736
rect 22560 16720 22612 16726
rect 22560 16662 22612 16668
rect 22744 16584 22796 16590
rect 22744 16526 22796 16532
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 22284 16040 22336 16046
rect 22756 16028 22784 16526
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 22836 16040 22888 16046
rect 22756 16000 22836 16028
rect 22284 15982 22336 15988
rect 22836 15982 22888 15988
rect 22192 15972 22244 15978
rect 22192 15914 22244 15920
rect 22296 15638 22324 15982
rect 22008 15632 22060 15638
rect 22008 15574 22060 15580
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22836 15564 22888 15570
rect 22836 15506 22888 15512
rect 22376 15496 22428 15502
rect 22376 15438 22428 15444
rect 22388 14958 22416 15438
rect 22744 15020 22796 15026
rect 22744 14962 22796 14968
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 21318 14716 21614 14736
rect 21374 14714 21398 14716
rect 21454 14714 21478 14716
rect 21534 14714 21558 14716
rect 21396 14662 21398 14714
rect 21460 14662 21472 14714
rect 21534 14662 21536 14714
rect 21374 14660 21398 14662
rect 21454 14660 21478 14662
rect 21534 14660 21558 14662
rect 21318 14640 21614 14660
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20168 14340 20220 14346
rect 20168 14282 20220 14288
rect 19800 13388 19852 13394
rect 19800 13330 19852 13336
rect 19708 12368 19760 12374
rect 19708 12310 19760 12316
rect 19812 12306 19840 13330
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 20088 11898 20116 12718
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19720 11218 19748 11630
rect 19904 11218 19932 11834
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19616 11144 19668 11150
rect 19616 11086 19668 11092
rect 19628 10674 19656 11086
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19616 10192 19668 10198
rect 19616 10134 19668 10140
rect 19628 9994 19656 10134
rect 19616 9988 19668 9994
rect 19616 9930 19668 9936
rect 19616 9648 19668 9654
rect 19614 9616 19616 9625
rect 19668 9616 19670 9625
rect 19524 9580 19576 9586
rect 19614 9551 19670 9560
rect 19524 9522 19576 9528
rect 19720 9518 19748 10542
rect 20180 10470 20208 14282
rect 20350 13152 20406 13161
rect 20350 13087 20406 13096
rect 20364 12986 20392 13087
rect 20442 13016 20498 13025
rect 20352 12980 20404 12986
rect 20442 12951 20498 12960
rect 20352 12922 20404 12928
rect 20456 12918 20484 12951
rect 20444 12912 20496 12918
rect 20444 12854 20496 12860
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20272 11762 20300 12718
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20272 11150 20300 11698
rect 20640 11558 20668 12786
rect 20732 11608 20760 14486
rect 22388 14414 22416 14894
rect 22376 14408 22428 14414
rect 22376 14350 22428 14356
rect 22376 14272 22428 14278
rect 22376 14214 22428 14220
rect 22388 13870 22416 14214
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 20904 13864 20956 13870
rect 22100 13864 22152 13870
rect 20904 13806 20956 13812
rect 22020 13812 22100 13818
rect 22020 13806 22152 13812
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22376 13864 22428 13870
rect 22376 13806 22428 13812
rect 20916 13462 20944 13806
rect 22020 13790 22140 13806
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21318 13628 21614 13648
rect 21374 13626 21398 13628
rect 21454 13626 21478 13628
rect 21534 13626 21558 13628
rect 21396 13574 21398 13626
rect 21460 13574 21472 13626
rect 21534 13574 21536 13626
rect 21374 13572 21398 13574
rect 21454 13572 21478 13574
rect 21534 13572 21558 13574
rect 21318 13552 21614 13572
rect 20904 13456 20956 13462
rect 20904 13398 20956 13404
rect 21744 13394 21772 13670
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 21732 13388 21784 13394
rect 21732 13330 21784 13336
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20824 11801 20852 12718
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 20810 11792 20866 11801
rect 21100 11762 21128 12174
rect 20810 11727 20812 11736
rect 20864 11727 20866 11736
rect 21088 11756 21140 11762
rect 20812 11698 20864 11704
rect 21088 11698 21140 11704
rect 20824 11667 20852 11698
rect 20904 11620 20956 11626
rect 20732 11580 20904 11608
rect 20904 11562 20956 11568
rect 20628 11552 20680 11558
rect 20628 11494 20680 11500
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 20628 11280 20680 11286
rect 21100 11257 21128 11290
rect 20628 11222 20680 11228
rect 21086 11248 21142 11257
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20640 10742 20668 11222
rect 21086 11183 21142 11192
rect 20904 11144 20956 11150
rect 20902 11112 20904 11121
rect 20956 11112 20958 11121
rect 20902 11047 20958 11056
rect 20902 10840 20958 10849
rect 20902 10775 20904 10784
rect 20956 10775 20958 10784
rect 20904 10746 20956 10752
rect 20628 10736 20680 10742
rect 20628 10678 20680 10684
rect 20812 10600 20864 10606
rect 20812 10542 20864 10548
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 20824 9761 20852 10542
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 20994 10024 21050 10033
rect 20994 9959 21050 9968
rect 20810 9752 20866 9761
rect 20810 9687 20866 9696
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 19708 9512 19760 9518
rect 19708 9454 19760 9460
rect 20732 9110 20760 9590
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20916 9110 20944 9454
rect 21008 9382 21036 9959
rect 21100 9450 21128 10066
rect 21192 9926 21220 13330
rect 21318 12540 21614 12560
rect 21374 12538 21398 12540
rect 21454 12538 21478 12540
rect 21534 12538 21558 12540
rect 21396 12486 21398 12538
rect 21460 12486 21472 12538
rect 21534 12486 21536 12538
rect 21374 12484 21398 12486
rect 21454 12484 21478 12486
rect 21534 12484 21558 12486
rect 21318 12464 21614 12484
rect 21640 12368 21692 12374
rect 21640 12310 21692 12316
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21560 11898 21588 12106
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21318 11452 21614 11472
rect 21374 11450 21398 11452
rect 21454 11450 21478 11452
rect 21534 11450 21558 11452
rect 21396 11398 21398 11450
rect 21460 11398 21472 11450
rect 21534 11398 21536 11450
rect 21374 11396 21398 11398
rect 21454 11396 21478 11398
rect 21534 11396 21558 11398
rect 21318 11376 21614 11396
rect 21652 11354 21680 12310
rect 21744 12306 21772 13330
rect 21732 12300 21784 12306
rect 21732 12242 21784 12248
rect 22020 12170 22048 13790
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22008 12164 22060 12170
rect 22008 12106 22060 12112
rect 22112 11898 22140 12718
rect 22296 12442 22324 13806
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21744 11082 21772 11698
rect 22480 11558 22508 14010
rect 22652 13524 22704 13530
rect 22652 13466 22704 13472
rect 22664 12889 22692 13466
rect 22650 12880 22706 12889
rect 22650 12815 22706 12824
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 21732 11076 21784 11082
rect 21732 11018 21784 11024
rect 22560 11008 22612 11014
rect 22560 10950 22612 10956
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 21318 10364 21614 10384
rect 21374 10362 21398 10364
rect 21454 10362 21478 10364
rect 21534 10362 21558 10364
rect 21396 10310 21398 10362
rect 21460 10310 21472 10362
rect 21534 10310 21536 10362
rect 21374 10308 21398 10310
rect 21454 10308 21478 10310
rect 21534 10308 21558 10310
rect 21318 10288 21614 10308
rect 22204 10130 22232 10610
rect 22572 10538 22600 10950
rect 22560 10532 22612 10538
rect 22560 10474 22612 10480
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 22192 10124 22244 10130
rect 22192 10066 22244 10072
rect 21284 9994 21312 10066
rect 21272 9988 21324 9994
rect 21272 9930 21324 9936
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 21088 9444 21140 9450
rect 21088 9386 21140 9392
rect 20996 9376 21048 9382
rect 21284 9364 21312 9930
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 20996 9318 21048 9324
rect 21192 9336 21312 9364
rect 21640 9376 21692 9382
rect 20720 9104 20772 9110
rect 20258 9072 20314 9081
rect 20720 9046 20772 9052
rect 20904 9104 20956 9110
rect 20904 9046 20956 9052
rect 20258 9007 20314 9016
rect 19616 8968 19668 8974
rect 19444 8928 19616 8956
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17972 5370 18000 5510
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 18236 5092 18288 5098
rect 18236 5034 18288 5040
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 17880 4622 17908 4966
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 18248 4554 18276 5034
rect 18236 4548 18288 4554
rect 18236 4490 18288 4496
rect 18234 4312 18290 4321
rect 18234 4247 18290 4256
rect 18248 4146 18276 4247
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18328 4004 18380 4010
rect 18328 3946 18380 3952
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 17788 3194 17816 3402
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 18248 3058 18276 3402
rect 18340 3058 18368 3946
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 17972 2310 18000 2790
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 18340 2106 18368 2382
rect 18328 2100 18380 2106
rect 18328 2042 18380 2048
rect 18524 800 18552 3470
rect 18708 2990 18736 6054
rect 19340 5772 19392 5778
rect 19260 5732 19340 5760
rect 18786 4584 18842 4593
rect 18786 4519 18842 4528
rect 18970 4584 19026 4593
rect 19260 4554 19288 5732
rect 19340 5714 19392 5720
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 18970 4519 19026 4528
rect 19248 4548 19300 4554
rect 18800 4078 18828 4519
rect 18984 4486 19012 4519
rect 19248 4490 19300 4496
rect 18880 4480 18932 4486
rect 18880 4422 18932 4428
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18892 3942 18920 4422
rect 19246 4312 19302 4321
rect 19352 4264 19380 5510
rect 19302 4256 19380 4264
rect 19246 4247 19380 4256
rect 19260 4236 19380 4247
rect 19338 4176 19394 4185
rect 19338 4111 19394 4120
rect 19064 4072 19116 4078
rect 18984 4032 19064 4060
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18800 2990 18828 3878
rect 18892 3602 18920 3878
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18708 2825 18736 2926
rect 18788 2848 18840 2854
rect 18694 2816 18750 2825
rect 18788 2790 18840 2796
rect 18694 2751 18750 2760
rect 18800 2689 18828 2790
rect 18786 2680 18842 2689
rect 18786 2615 18842 2624
rect 18984 1970 19012 4032
rect 19248 4072 19300 4078
rect 19064 4014 19116 4020
rect 19168 4020 19248 4026
rect 19168 4014 19300 4020
rect 19168 3998 19288 4014
rect 19168 3913 19196 3998
rect 19154 3904 19210 3913
rect 19154 3839 19210 3848
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 19076 2990 19104 3674
rect 19352 3602 19380 4111
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 19260 2990 19288 3538
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 18972 1964 19024 1970
rect 18972 1906 19024 1912
rect 19444 800 19472 8570
rect 19536 7954 19564 8928
rect 19616 8910 19668 8916
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 19800 8832 19852 8838
rect 20088 8786 20116 8910
rect 19852 8780 20116 8786
rect 19800 8774 20116 8780
rect 19812 8758 20116 8774
rect 20088 8430 20116 8758
rect 20166 8528 20222 8537
rect 20166 8463 20168 8472
rect 20220 8463 20222 8472
rect 20168 8434 20220 8440
rect 20076 8424 20128 8430
rect 20076 8366 20128 8372
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19536 7546 19564 7890
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19720 7206 19748 8026
rect 19996 7546 20024 8230
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 20088 7410 20116 8230
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 19708 7200 19760 7206
rect 19708 7142 19760 7148
rect 19720 6866 19748 7142
rect 20272 6934 20300 9007
rect 21192 8974 21220 9336
rect 21640 9318 21692 9324
rect 21318 9276 21614 9296
rect 21374 9274 21398 9276
rect 21454 9274 21478 9276
rect 21534 9274 21558 9276
rect 21396 9222 21398 9274
rect 21460 9222 21472 9274
rect 21534 9222 21536 9274
rect 21374 9220 21398 9222
rect 21454 9220 21478 9222
rect 21534 9220 21558 9222
rect 21318 9200 21614 9220
rect 21546 9072 21602 9081
rect 21546 9007 21548 9016
rect 21600 9007 21602 9016
rect 21548 8978 21600 8984
rect 21180 8968 21232 8974
rect 20902 8936 20958 8945
rect 21180 8910 21232 8916
rect 20902 8871 20958 8880
rect 20916 8838 20944 8871
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20718 8664 20774 8673
rect 20718 8599 20774 8608
rect 20732 8566 20760 8599
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20824 8430 20852 8774
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 20548 8022 20576 8366
rect 20444 8016 20496 8022
rect 20444 7958 20496 7964
rect 20536 8016 20588 8022
rect 20536 7958 20588 7964
rect 20456 7857 20484 7958
rect 20548 7886 20576 7958
rect 20640 7954 20668 8366
rect 20824 7954 20852 8366
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20812 7948 20864 7954
rect 20812 7890 20864 7896
rect 20536 7880 20588 7886
rect 20442 7848 20498 7857
rect 20536 7822 20588 7828
rect 20442 7783 20498 7792
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20364 7478 20392 7686
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 20640 7410 20668 7890
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20260 6928 20312 6934
rect 20260 6870 20312 6876
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19536 6322 19564 6734
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20074 6488 20130 6497
rect 20074 6423 20130 6432
rect 20088 6390 20116 6423
rect 19892 6384 19944 6390
rect 19892 6326 19944 6332
rect 20076 6384 20128 6390
rect 20076 6326 20128 6332
rect 20168 6384 20220 6390
rect 20168 6326 20220 6332
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19904 5166 19932 6326
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 20088 5234 20116 5646
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 19892 5160 19944 5166
rect 19892 5102 19944 5108
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19996 4214 20024 5102
rect 19984 4208 20036 4214
rect 19984 4150 20036 4156
rect 20180 4146 20208 6326
rect 20272 6254 20300 6598
rect 20350 6352 20406 6361
rect 20732 6322 20760 7822
rect 20350 6287 20406 6296
rect 20720 6316 20772 6322
rect 20364 6254 20392 6287
rect 20720 6258 20772 6264
rect 20824 6254 20852 7890
rect 20916 7274 20944 8298
rect 21318 8188 21614 8208
rect 21374 8186 21398 8188
rect 21454 8186 21478 8188
rect 21534 8186 21558 8188
rect 21396 8134 21398 8186
rect 21460 8134 21472 8186
rect 21534 8134 21536 8186
rect 21374 8132 21398 8134
rect 21454 8132 21478 8134
rect 21534 8132 21558 8134
rect 21318 8112 21614 8132
rect 21088 7948 21140 7954
rect 21088 7890 21140 7896
rect 20904 7268 20956 7274
rect 20904 7210 20956 7216
rect 20916 6866 20944 7210
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 21008 6769 21036 6802
rect 20994 6760 21050 6769
rect 20994 6695 21050 6704
rect 20260 6248 20312 6254
rect 20260 6190 20312 6196
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 20088 3942 20116 4014
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19720 2446 19748 3334
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 20272 800 20300 6190
rect 20364 4486 20392 6190
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20534 4040 20590 4049
rect 20364 3398 20392 4014
rect 20534 3975 20590 3984
rect 20548 3942 20576 3975
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20640 3466 20668 5170
rect 20812 4004 20864 4010
rect 20812 3946 20864 3952
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 20352 3392 20404 3398
rect 20352 3334 20404 3340
rect 20640 2990 20668 3402
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20732 2446 20760 3470
rect 20824 2990 20852 3946
rect 20916 3602 20944 5306
rect 21008 4690 21036 6695
rect 21100 5778 21128 7890
rect 21318 7100 21614 7120
rect 21374 7098 21398 7100
rect 21454 7098 21478 7100
rect 21534 7098 21558 7100
rect 21396 7046 21398 7098
rect 21460 7046 21472 7098
rect 21534 7046 21536 7098
rect 21374 7044 21398 7046
rect 21454 7044 21478 7046
rect 21534 7044 21558 7046
rect 21318 7024 21614 7044
rect 21652 6916 21680 9318
rect 21744 9194 21772 9454
rect 21836 9330 21864 10066
rect 22192 9512 22244 9518
rect 22192 9454 22244 9460
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 21836 9302 21956 9330
rect 21744 9166 21864 9194
rect 21836 9110 21864 9166
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 21836 8634 21864 8910
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21822 8392 21878 8401
rect 21822 8327 21824 8336
rect 21876 8327 21878 8336
rect 21928 8344 21956 9302
rect 22020 8956 22048 9386
rect 22100 8968 22152 8974
rect 22020 8928 22100 8956
rect 22100 8910 22152 8916
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 22020 8537 22048 8570
rect 22204 8566 22232 9454
rect 22284 9036 22336 9042
rect 22336 8996 22508 9024
rect 22284 8978 22336 8984
rect 22376 8900 22428 8906
rect 22376 8842 22428 8848
rect 22388 8566 22416 8842
rect 22192 8560 22244 8566
rect 22006 8528 22062 8537
rect 22192 8502 22244 8508
rect 22376 8560 22428 8566
rect 22376 8502 22428 8508
rect 22006 8463 22062 8472
rect 22204 8430 22232 8502
rect 22480 8498 22508 8996
rect 22560 8900 22612 8906
rect 22560 8842 22612 8848
rect 22572 8673 22600 8842
rect 22558 8664 22614 8673
rect 22558 8599 22614 8608
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 21928 8316 22048 8344
rect 21824 8298 21876 8304
rect 21560 6888 21680 6916
rect 21560 6254 21588 6888
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 21730 6216 21786 6225
rect 21730 6151 21786 6160
rect 21744 6118 21772 6151
rect 21732 6112 21784 6118
rect 21732 6054 21784 6060
rect 21318 6012 21614 6032
rect 21374 6010 21398 6012
rect 21454 6010 21478 6012
rect 21534 6010 21558 6012
rect 21396 5958 21398 6010
rect 21460 5958 21472 6010
rect 21534 5958 21536 6010
rect 21374 5956 21398 5958
rect 21454 5956 21478 5958
rect 21534 5956 21558 5958
rect 21318 5936 21614 5956
rect 21180 5840 21232 5846
rect 21180 5782 21232 5788
rect 21088 5772 21140 5778
rect 21088 5714 21140 5720
rect 21192 5545 21220 5782
rect 21178 5536 21234 5545
rect 21178 5471 21234 5480
rect 21192 5098 21220 5471
rect 21180 5092 21232 5098
rect 21180 5034 21232 5040
rect 21318 4924 21614 4944
rect 21374 4922 21398 4924
rect 21454 4922 21478 4924
rect 21534 4922 21558 4924
rect 21396 4870 21398 4922
rect 21460 4870 21472 4922
rect 21534 4870 21536 4922
rect 21374 4868 21398 4870
rect 21454 4868 21478 4870
rect 21534 4868 21558 4870
rect 21318 4848 21614 4868
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 21318 3836 21614 3856
rect 21374 3834 21398 3836
rect 21454 3834 21478 3836
rect 21534 3834 21558 3836
rect 21396 3782 21398 3834
rect 21460 3782 21472 3834
rect 21534 3782 21536 3834
rect 21374 3780 21398 3782
rect 21454 3780 21478 3782
rect 21534 3780 21558 3782
rect 21318 3760 21614 3780
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 20824 2582 20852 2926
rect 20812 2576 20864 2582
rect 20812 2518 20864 2524
rect 21100 2514 21128 3674
rect 21180 3188 21232 3194
rect 21180 3130 21232 3136
rect 21088 2508 21140 2514
rect 21088 2450 21140 2456
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 21192 800 21220 3130
rect 21836 3058 21864 8298
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 21928 6254 21956 7346
rect 22020 7342 22048 8316
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 22112 7886 22140 8026
rect 22204 7954 22232 8026
rect 22192 7948 22244 7954
rect 22192 7890 22244 7896
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 22284 7880 22336 7886
rect 22284 7822 22336 7828
rect 22296 7478 22324 7822
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 22480 7274 22508 7754
rect 22468 7268 22520 7274
rect 22468 7210 22520 7216
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 21928 4622 21956 6190
rect 22388 5642 22416 6734
rect 22376 5636 22428 5642
rect 22376 5578 22428 5584
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 22006 3360 22062 3369
rect 22006 3295 22062 3304
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21318 2748 21614 2768
rect 21374 2746 21398 2748
rect 21454 2746 21478 2748
rect 21534 2746 21558 2748
rect 21396 2694 21398 2746
rect 21460 2694 21472 2746
rect 21534 2694 21536 2746
rect 21374 2692 21398 2694
rect 21454 2692 21478 2694
rect 21534 2692 21558 2694
rect 21318 2672 21614 2692
rect 21732 2304 21784 2310
rect 21732 2246 21784 2252
rect 21744 2106 21772 2246
rect 21732 2100 21784 2106
rect 21732 2042 21784 2048
rect 22020 800 22048 3295
rect 22388 2961 22416 5578
rect 22468 4684 22520 4690
rect 22468 4626 22520 4632
rect 22480 4282 22508 4626
rect 22572 4622 22600 7890
rect 22664 7857 22692 11154
rect 22756 8906 22784 14962
rect 22848 13190 22876 15506
rect 22940 14822 22968 16390
rect 23032 15162 23060 16526
rect 23664 16244 23716 16250
rect 23664 16186 23716 16192
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 23020 15156 23072 15162
rect 23020 15098 23072 15104
rect 23020 14952 23072 14958
rect 23020 14894 23072 14900
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 23032 14346 23060 14894
rect 23020 14340 23072 14346
rect 23020 14282 23072 14288
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 23032 13433 23060 13874
rect 23018 13424 23074 13433
rect 23018 13359 23020 13368
rect 23072 13359 23074 13368
rect 23020 13330 23072 13336
rect 22836 13184 22888 13190
rect 22836 13126 22888 13132
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22744 8900 22796 8906
rect 22744 8842 22796 8848
rect 22940 7886 22968 9862
rect 23124 9654 23152 15506
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 23308 14958 23336 15438
rect 23676 15434 23704 16186
rect 24044 16046 24072 17070
rect 24032 16040 24084 16046
rect 24084 16000 24164 16028
rect 24032 15982 24084 15988
rect 23664 15428 23716 15434
rect 23664 15370 23716 15376
rect 23676 15026 23704 15370
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23492 11694 23520 12174
rect 23584 12102 23612 12242
rect 23676 12102 23704 12718
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23664 12096 23716 12102
rect 23664 12038 23716 12044
rect 23756 11824 23808 11830
rect 23754 11792 23756 11801
rect 23808 11792 23810 11801
rect 23754 11727 23810 11736
rect 23480 11688 23532 11694
rect 23480 11630 23532 11636
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 23308 9994 23336 11154
rect 23388 11008 23440 11014
rect 23388 10950 23440 10956
rect 23400 10130 23428 10950
rect 23572 10600 23624 10606
rect 23572 10542 23624 10548
rect 23584 10130 23612 10542
rect 23860 10470 23888 12378
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 23296 9988 23348 9994
rect 23296 9930 23348 9936
rect 23112 9648 23164 9654
rect 23756 9648 23808 9654
rect 23112 9590 23164 9596
rect 23754 9616 23756 9625
rect 23808 9616 23810 9625
rect 23124 9042 23152 9590
rect 23952 9586 23980 12718
rect 24044 11694 24072 14758
rect 24136 14006 24164 16000
rect 24860 15972 24912 15978
rect 24860 15914 24912 15920
rect 24492 15564 24544 15570
rect 24492 15506 24544 15512
rect 24504 14550 24532 15506
rect 24872 14618 24900 15914
rect 24964 15638 24992 17070
rect 24952 15632 25004 15638
rect 24952 15574 25004 15580
rect 25424 14958 25452 17274
rect 25884 17202 25912 18835
rect 27724 17338 27752 18835
rect 27712 17332 27764 17338
rect 27712 17274 27764 17280
rect 25872 17196 25924 17202
rect 25872 17138 25924 17144
rect 25884 16250 25912 17138
rect 29656 17134 29684 18835
rect 31588 17626 31616 18835
rect 31404 17598 31616 17626
rect 29644 17128 29696 17134
rect 29644 17070 29696 17076
rect 27252 17060 27304 17066
rect 27252 17002 27304 17008
rect 25872 16244 25924 16250
rect 25872 16186 25924 16192
rect 27068 15904 27120 15910
rect 27068 15846 27120 15852
rect 27080 15706 27108 15846
rect 27068 15700 27120 15706
rect 27068 15642 27120 15648
rect 27080 15570 27108 15642
rect 27068 15564 27120 15570
rect 27068 15506 27120 15512
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 25516 15162 25544 15438
rect 27264 15434 27292 17002
rect 28172 16992 28224 16998
rect 28172 16934 28224 16940
rect 27988 16584 28040 16590
rect 27988 16526 28040 16532
rect 27896 16176 27948 16182
rect 27896 16118 27948 16124
rect 27528 15564 27580 15570
rect 27528 15506 27580 15512
rect 27252 15428 27304 15434
rect 27252 15370 27304 15376
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 25412 14952 25464 14958
rect 25412 14894 25464 14900
rect 25504 14952 25556 14958
rect 25504 14894 25556 14900
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24492 14544 24544 14550
rect 24492 14486 24544 14492
rect 24308 14476 24360 14482
rect 24308 14418 24360 14424
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24320 14074 24348 14418
rect 24308 14068 24360 14074
rect 24308 14010 24360 14016
rect 24124 14000 24176 14006
rect 24124 13942 24176 13948
rect 24400 13524 24452 13530
rect 24400 13466 24452 13472
rect 24216 13388 24268 13394
rect 24216 13330 24268 13336
rect 24124 12300 24176 12306
rect 24124 12242 24176 12248
rect 24032 11688 24084 11694
rect 24032 11630 24084 11636
rect 24136 9654 24164 12242
rect 24228 11218 24256 13330
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 24320 12986 24348 13126
rect 24308 12980 24360 12986
rect 24308 12922 24360 12928
rect 24320 12238 24348 12922
rect 24412 12646 24440 13466
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 24412 12442 24440 12582
rect 24400 12436 24452 12442
rect 24400 12378 24452 12384
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 24216 11212 24268 11218
rect 24216 11154 24268 11160
rect 24228 10674 24256 11154
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24124 9648 24176 9654
rect 24124 9590 24176 9596
rect 23754 9551 23810 9560
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 24228 9518 24256 10610
rect 24688 10062 24716 14418
rect 25228 13388 25280 13394
rect 25228 13330 25280 13336
rect 25240 12306 25268 13330
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 25412 12300 25464 12306
rect 25516 12288 25544 14894
rect 27264 14890 27292 15370
rect 27540 15366 27568 15506
rect 27908 15434 27936 16118
rect 28000 16114 28028 16526
rect 27988 16108 28040 16114
rect 27988 16050 28040 16056
rect 28184 15978 28212 16934
rect 29656 16726 29684 17070
rect 30196 17060 30248 17066
rect 30196 17002 30248 17008
rect 30208 16726 30236 17002
rect 29644 16720 29696 16726
rect 29644 16662 29696 16668
rect 30196 16720 30248 16726
rect 30196 16662 30248 16668
rect 31404 16658 31432 17598
rect 31500 17436 31796 17456
rect 31556 17434 31580 17436
rect 31636 17434 31660 17436
rect 31716 17434 31740 17436
rect 31578 17382 31580 17434
rect 31642 17382 31654 17434
rect 31716 17382 31718 17434
rect 31556 17380 31580 17382
rect 31636 17380 31660 17382
rect 31716 17380 31740 17382
rect 31500 17360 31796 17380
rect 33520 17134 33548 18835
rect 33508 17128 33560 17134
rect 33508 17070 33560 17076
rect 33520 16794 33548 17070
rect 34244 16992 34296 16998
rect 34244 16934 34296 16940
rect 34888 16992 34940 16998
rect 34888 16934 34940 16940
rect 33508 16788 33560 16794
rect 33508 16730 33560 16736
rect 29276 16652 29328 16658
rect 29276 16594 29328 16600
rect 31392 16652 31444 16658
rect 31392 16594 31444 16600
rect 28724 16448 28776 16454
rect 28724 16390 28776 16396
rect 28172 15972 28224 15978
rect 28172 15914 28224 15920
rect 28736 15638 28764 16390
rect 29288 16046 29316 16594
rect 31404 16250 31432 16594
rect 32864 16584 32916 16590
rect 32864 16526 32916 16532
rect 31500 16348 31796 16368
rect 31556 16346 31580 16348
rect 31636 16346 31660 16348
rect 31716 16346 31740 16348
rect 31578 16294 31580 16346
rect 31642 16294 31654 16346
rect 31716 16294 31718 16346
rect 31556 16292 31580 16294
rect 31636 16292 31660 16294
rect 31716 16292 31740 16294
rect 31500 16272 31796 16292
rect 31392 16244 31444 16250
rect 31392 16186 31444 16192
rect 29276 16040 29328 16046
rect 29276 15982 29328 15988
rect 29552 16040 29604 16046
rect 29552 15982 29604 15988
rect 28724 15632 28776 15638
rect 28724 15574 28776 15580
rect 28632 15564 28684 15570
rect 28632 15506 28684 15512
rect 28816 15564 28868 15570
rect 28868 15524 28948 15552
rect 28816 15506 28868 15512
rect 27896 15428 27948 15434
rect 27896 15370 27948 15376
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27908 15162 27936 15370
rect 28644 15162 28672 15506
rect 27896 15156 27948 15162
rect 27896 15098 27948 15104
rect 28632 15156 28684 15162
rect 28632 15098 28684 15104
rect 28172 15088 28224 15094
rect 28172 15030 28224 15036
rect 27896 14952 27948 14958
rect 27896 14894 27948 14900
rect 27252 14884 27304 14890
rect 27252 14826 27304 14832
rect 27908 14482 27936 14894
rect 26608 14476 26660 14482
rect 26608 14418 26660 14424
rect 26792 14476 26844 14482
rect 26792 14418 26844 14424
rect 27896 14476 27948 14482
rect 27896 14418 27948 14424
rect 26620 13938 26648 14418
rect 25872 13932 25924 13938
rect 25872 13874 25924 13880
rect 26608 13932 26660 13938
rect 26608 13874 26660 13880
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25792 12918 25820 13126
rect 25780 12912 25832 12918
rect 25780 12854 25832 12860
rect 25464 12260 25544 12288
rect 25412 12242 25464 12248
rect 24952 12164 25004 12170
rect 24952 12106 25004 12112
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24780 10674 24808 11630
rect 24964 11121 24992 12106
rect 24950 11112 25006 11121
rect 24950 11047 25006 11056
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24780 10198 24808 10610
rect 24768 10192 24820 10198
rect 24768 10134 24820 10140
rect 24676 10056 24728 10062
rect 24676 9998 24728 10004
rect 23204 9512 23256 9518
rect 23204 9454 23256 9460
rect 24216 9512 24268 9518
rect 24216 9454 24268 9460
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23216 8906 23244 9454
rect 24780 9042 24808 10134
rect 24964 9110 24992 11047
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 25056 9926 25084 10066
rect 25044 9920 25096 9926
rect 25044 9862 25096 9868
rect 25240 9625 25268 12242
rect 25320 11552 25372 11558
rect 25320 11494 25372 11500
rect 25332 10062 25360 11494
rect 25424 10606 25452 12242
rect 25504 12096 25556 12102
rect 25504 12038 25556 12044
rect 25516 11898 25544 12038
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 25780 11688 25832 11694
rect 25780 11630 25832 11636
rect 25412 10600 25464 10606
rect 25412 10542 25464 10548
rect 25792 10538 25820 11630
rect 25884 10674 25912 13874
rect 26148 13864 26200 13870
rect 26148 13806 26200 13812
rect 26160 12918 26188 13806
rect 26240 13252 26292 13258
rect 26240 13194 26292 13200
rect 26252 12918 26280 13194
rect 26148 12912 26200 12918
rect 26148 12854 26200 12860
rect 26240 12912 26292 12918
rect 26240 12854 26292 12860
rect 26620 12850 26648 13874
rect 26804 13530 26832 14418
rect 27068 13796 27120 13802
rect 27068 13738 27120 13744
rect 26792 13524 26844 13530
rect 26792 13466 26844 13472
rect 26884 13524 26936 13530
rect 26884 13466 26936 13472
rect 26896 13025 26924 13466
rect 27080 13394 27108 13738
rect 27068 13388 27120 13394
rect 27068 13330 27120 13336
rect 27344 13388 27396 13394
rect 27344 13330 27396 13336
rect 27988 13388 28040 13394
rect 27988 13330 28040 13336
rect 27080 13161 27108 13330
rect 27066 13152 27122 13161
rect 27066 13087 27122 13096
rect 26882 13016 26938 13025
rect 26882 12951 26938 12960
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 26792 12776 26844 12782
rect 26792 12718 26844 12724
rect 26332 12708 26384 12714
rect 26332 12650 26384 12656
rect 26344 12617 26372 12650
rect 26330 12608 26386 12617
rect 26330 12543 26386 12552
rect 26804 11694 26832 12718
rect 27356 11762 27384 13330
rect 27710 12880 27766 12889
rect 27710 12815 27766 12824
rect 27724 12782 27752 12815
rect 27712 12776 27764 12782
rect 27712 12718 27764 12724
rect 27620 12640 27672 12646
rect 27896 12640 27948 12646
rect 27620 12582 27672 12588
rect 27894 12608 27896 12617
rect 27948 12608 27950 12617
rect 27632 11762 27660 12582
rect 27894 12543 27950 12552
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27620 11756 27672 11762
rect 27620 11698 27672 11704
rect 27896 11756 27948 11762
rect 27896 11698 27948 11704
rect 26148 11688 26200 11694
rect 26148 11630 26200 11636
rect 26792 11688 26844 11694
rect 27804 11688 27856 11694
rect 26792 11630 26844 11636
rect 27356 11636 27804 11642
rect 27356 11630 27856 11636
rect 26056 11552 26108 11558
rect 26056 11494 26108 11500
rect 26068 11218 26096 11494
rect 26056 11212 26108 11218
rect 26056 11154 26108 11160
rect 25872 10668 25924 10674
rect 25872 10610 25924 10616
rect 25780 10532 25832 10538
rect 25780 10474 25832 10480
rect 25792 10198 25820 10474
rect 26160 10470 26188 11630
rect 27356 11626 27844 11630
rect 27344 11620 27844 11626
rect 27396 11614 27844 11620
rect 27344 11562 27396 11568
rect 27160 11280 27212 11286
rect 27160 11222 27212 11228
rect 26700 11008 26752 11014
rect 26700 10950 26752 10956
rect 27068 11008 27120 11014
rect 27068 10950 27120 10956
rect 26148 10464 26200 10470
rect 26148 10406 26200 10412
rect 25780 10192 25832 10198
rect 25780 10134 25832 10140
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25226 9616 25282 9625
rect 25226 9551 25282 9560
rect 25332 9518 25360 9998
rect 26160 9586 26188 10406
rect 26424 10124 26476 10130
rect 26424 10066 26476 10072
rect 26436 9586 26464 10066
rect 26712 9994 26740 10950
rect 27080 10674 27108 10950
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 27172 10554 27200 11222
rect 27080 10526 27200 10554
rect 26884 10464 26936 10470
rect 26884 10406 26936 10412
rect 26896 10130 26924 10406
rect 27080 10130 27108 10526
rect 27540 10470 27568 11614
rect 27802 11248 27858 11257
rect 27620 11212 27672 11218
rect 27908 11218 27936 11698
rect 28000 11558 28028 13330
rect 28080 12232 28132 12238
rect 28080 12174 28132 12180
rect 28092 11762 28120 12174
rect 28080 11756 28132 11762
rect 28080 11698 28132 11704
rect 27988 11552 28040 11558
rect 27988 11494 28040 11500
rect 27802 11183 27858 11192
rect 27896 11212 27948 11218
rect 27620 11154 27672 11160
rect 27632 10674 27660 11154
rect 27816 11150 27844 11183
rect 27896 11154 27948 11160
rect 27804 11144 27856 11150
rect 27804 11086 27856 11092
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 27620 10532 27672 10538
rect 27620 10474 27672 10480
rect 27528 10464 27580 10470
rect 27528 10406 27580 10412
rect 27632 10130 27660 10474
rect 26884 10124 26936 10130
rect 26884 10066 26936 10072
rect 27068 10124 27120 10130
rect 27068 10066 27120 10072
rect 27620 10124 27672 10130
rect 27620 10066 27672 10072
rect 26700 9988 26752 9994
rect 26700 9930 26752 9936
rect 26148 9580 26200 9586
rect 26148 9522 26200 9528
rect 26424 9580 26476 9586
rect 26424 9522 26476 9528
rect 25320 9512 25372 9518
rect 25320 9454 25372 9460
rect 27080 9450 27108 10066
rect 27436 9988 27488 9994
rect 27436 9930 27488 9936
rect 27712 9988 27764 9994
rect 27712 9930 27764 9936
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 26516 9444 26568 9450
rect 26516 9386 26568 9392
rect 27068 9444 27120 9450
rect 27068 9386 27120 9392
rect 24952 9104 25004 9110
rect 24952 9046 25004 9052
rect 24768 9036 24820 9042
rect 24768 8978 24820 8984
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 24952 8968 25004 8974
rect 24952 8910 25004 8916
rect 23204 8900 23256 8906
rect 23204 8842 23256 8848
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 23400 8430 23428 8774
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 22928 7880 22980 7886
rect 22650 7848 22706 7857
rect 22928 7822 22980 7828
rect 22650 7783 22706 7792
rect 23296 7268 23348 7274
rect 23296 7210 23348 7216
rect 22744 6180 22796 6186
rect 22744 6122 22796 6128
rect 22756 4690 22784 6122
rect 23204 5908 23256 5914
rect 23204 5850 23256 5856
rect 23112 5568 23164 5574
rect 23112 5510 23164 5516
rect 23124 5370 23152 5510
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 23124 4758 23152 5306
rect 23112 4752 23164 4758
rect 23112 4694 23164 4700
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22468 4276 22520 4282
rect 22468 4218 22520 4224
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22468 3392 22520 3398
rect 22468 3334 22520 3340
rect 22480 3194 22508 3334
rect 22468 3188 22520 3194
rect 22468 3130 22520 3136
rect 22572 3097 22600 4082
rect 22926 4040 22982 4049
rect 22926 3975 22982 3984
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22664 3670 22692 3878
rect 22652 3664 22704 3670
rect 22652 3606 22704 3612
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 22558 3088 22614 3097
rect 22558 3023 22614 3032
rect 22572 2990 22600 3023
rect 22560 2984 22612 2990
rect 22374 2952 22430 2961
rect 22560 2926 22612 2932
rect 22374 2887 22430 2896
rect 22848 2854 22876 3470
rect 22836 2848 22888 2854
rect 22836 2790 22888 2796
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 22112 2106 22140 2586
rect 22848 2514 22876 2790
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 22100 2100 22152 2106
rect 22100 2042 22152 2048
rect 22940 800 22968 3975
rect 23216 3602 23244 5850
rect 23308 4010 23336 7210
rect 23400 6866 23428 8366
rect 23676 7954 23704 8910
rect 23848 8900 23900 8906
rect 23848 8842 23900 8848
rect 23860 8566 23888 8842
rect 23848 8560 23900 8566
rect 23848 8502 23900 8508
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 24216 7336 24268 7342
rect 24216 7278 24268 7284
rect 23388 6860 23440 6866
rect 23388 6802 23440 6808
rect 23572 6860 23624 6866
rect 23572 6802 23624 6808
rect 23584 6458 23612 6802
rect 23848 6792 23900 6798
rect 23848 6734 23900 6740
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 23480 5840 23532 5846
rect 23480 5782 23532 5788
rect 23296 4004 23348 4010
rect 23296 3946 23348 3952
rect 23492 3738 23520 5782
rect 23860 5574 23888 6734
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 23572 5568 23624 5574
rect 23572 5510 23624 5516
rect 23848 5568 23900 5574
rect 23848 5510 23900 5516
rect 23584 5302 23612 5510
rect 23572 5296 23624 5302
rect 23572 5238 23624 5244
rect 23664 5092 23716 5098
rect 23664 5034 23716 5040
rect 23676 4078 23704 5034
rect 23860 4078 23888 5510
rect 24044 5273 24072 6054
rect 24030 5264 24086 5273
rect 23952 5222 24030 5250
rect 23952 4185 23980 5222
rect 24030 5199 24086 5208
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 24044 4554 24072 5102
rect 24032 4548 24084 4554
rect 24032 4490 24084 4496
rect 23938 4176 23994 4185
rect 23938 4111 23994 4120
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 23848 4072 23900 4078
rect 23848 4014 23900 4020
rect 23480 3732 23532 3738
rect 23480 3674 23532 3680
rect 23204 3596 23256 3602
rect 23204 3538 23256 3544
rect 23676 3194 23704 4014
rect 24228 3602 24256 7278
rect 24872 5778 24900 8366
rect 24964 6254 24992 8910
rect 25412 8832 25464 8838
rect 25412 8774 25464 8780
rect 25424 8430 25452 8774
rect 26528 8498 26556 9386
rect 26608 8832 26660 8838
rect 26608 8774 26660 8780
rect 26516 8492 26568 8498
rect 26516 8434 26568 8440
rect 25412 8424 25464 8430
rect 25412 8366 25464 8372
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25780 7744 25832 7750
rect 25780 7686 25832 7692
rect 25044 7268 25096 7274
rect 25044 7210 25096 7216
rect 25056 6866 25084 7210
rect 25596 7200 25648 7206
rect 25596 7142 25648 7148
rect 25044 6860 25096 6866
rect 25044 6802 25096 6808
rect 25228 6724 25280 6730
rect 25228 6666 25280 6672
rect 25240 6322 25268 6666
rect 25228 6316 25280 6322
rect 25228 6258 25280 6264
rect 24952 6248 25004 6254
rect 24952 6190 25004 6196
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24320 4622 24348 5170
rect 24860 4684 24912 4690
rect 24860 4626 24912 4632
rect 24308 4616 24360 4622
rect 24308 4558 24360 4564
rect 24872 4146 24900 4626
rect 24860 4140 24912 4146
rect 24860 4082 24912 4088
rect 24582 3768 24638 3777
rect 24582 3703 24638 3712
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 23754 3224 23810 3233
rect 23664 3188 23716 3194
rect 23754 3159 23810 3168
rect 23664 3130 23716 3136
rect 23768 800 23796 3159
rect 24124 3120 24176 3126
rect 24124 3062 24176 3068
rect 24136 2689 24164 3062
rect 24308 2984 24360 2990
rect 24308 2926 24360 2932
rect 24122 2680 24178 2689
rect 24122 2615 24178 2624
rect 24320 2446 24348 2926
rect 24308 2440 24360 2446
rect 24308 2382 24360 2388
rect 24596 800 24624 3703
rect 24860 3528 24912 3534
rect 24860 3470 24912 3476
rect 24872 3058 24900 3470
rect 24860 3052 24912 3058
rect 24860 2994 24912 3000
rect 24964 2310 24992 6190
rect 25608 5846 25636 7142
rect 25700 6934 25728 7686
rect 25792 7478 25820 7686
rect 25780 7472 25832 7478
rect 25780 7414 25832 7420
rect 25688 6928 25740 6934
rect 25688 6870 25740 6876
rect 25964 6792 26016 6798
rect 25964 6734 26016 6740
rect 25976 6118 26004 6734
rect 26620 6662 26648 8774
rect 26884 8424 26936 8430
rect 27068 8424 27120 8430
rect 26936 8372 27068 8378
rect 27172 8401 27200 9522
rect 27252 9512 27304 9518
rect 27252 9454 27304 9460
rect 26884 8366 27120 8372
rect 27158 8392 27214 8401
rect 26896 8350 27108 8366
rect 27158 8327 27214 8336
rect 27160 7948 27212 7954
rect 27160 7890 27212 7896
rect 27172 7342 27200 7890
rect 27160 7336 27212 7342
rect 27160 7278 27212 7284
rect 27172 6934 27200 7278
rect 27160 6928 27212 6934
rect 27160 6870 27212 6876
rect 26884 6860 26936 6866
rect 26884 6802 26936 6808
rect 26976 6860 27028 6866
rect 26976 6802 27028 6808
rect 26608 6656 26660 6662
rect 26608 6598 26660 6604
rect 25964 6112 26016 6118
rect 25964 6054 26016 6060
rect 25596 5840 25648 5846
rect 25596 5782 25648 5788
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 25320 5772 25372 5778
rect 25320 5714 25372 5720
rect 25240 4826 25268 5714
rect 25332 5166 25360 5714
rect 26424 5636 26476 5642
rect 26424 5578 26476 5584
rect 25504 5364 25556 5370
rect 25504 5306 25556 5312
rect 25516 5166 25544 5306
rect 25320 5160 25372 5166
rect 25504 5160 25556 5166
rect 25320 5102 25372 5108
rect 25502 5128 25504 5137
rect 25964 5160 26016 5166
rect 25556 5128 25558 5137
rect 25964 5102 26016 5108
rect 25502 5063 25558 5072
rect 25228 4820 25280 4826
rect 25228 4762 25280 4768
rect 25412 4684 25464 4690
rect 25516 4672 25544 5063
rect 25976 5030 26004 5102
rect 25964 5024 26016 5030
rect 25964 4966 26016 4972
rect 26436 4690 26464 5578
rect 26620 5166 26648 6598
rect 26896 5302 26924 6802
rect 26988 5778 27016 6802
rect 27158 5944 27214 5953
rect 27264 5914 27292 9454
rect 27448 8974 27476 9930
rect 27620 9920 27672 9926
rect 27620 9862 27672 9868
rect 27528 9512 27580 9518
rect 27632 9500 27660 9862
rect 27580 9472 27660 9500
rect 27528 9454 27580 9460
rect 27724 9081 27752 9930
rect 27896 9648 27948 9654
rect 27896 9590 27948 9596
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27710 9072 27766 9081
rect 27816 9042 27844 9318
rect 27710 9007 27766 9016
rect 27804 9036 27856 9042
rect 27344 8968 27396 8974
rect 27344 8910 27396 8916
rect 27436 8968 27488 8974
rect 27436 8910 27488 8916
rect 27356 8022 27384 8910
rect 27436 8356 27488 8362
rect 27436 8298 27488 8304
rect 27620 8356 27672 8362
rect 27620 8298 27672 8304
rect 27344 8016 27396 8022
rect 27344 7958 27396 7964
rect 27448 7342 27476 8298
rect 27632 8022 27660 8298
rect 27620 8016 27672 8022
rect 27620 7958 27672 7964
rect 27724 7954 27752 9007
rect 27804 8978 27856 8984
rect 27816 8498 27844 8978
rect 27804 8492 27856 8498
rect 27804 8434 27856 8440
rect 27816 7954 27844 8434
rect 27712 7948 27764 7954
rect 27712 7890 27764 7896
rect 27804 7948 27856 7954
rect 27804 7890 27856 7896
rect 27908 7886 27936 9590
rect 27988 7948 28040 7954
rect 27988 7890 28040 7896
rect 27896 7880 27948 7886
rect 27896 7822 27948 7828
rect 28000 7478 28028 7890
rect 27988 7472 28040 7478
rect 27988 7414 28040 7420
rect 27436 7336 27488 7342
rect 27436 7278 27488 7284
rect 28078 7032 28134 7041
rect 28078 6967 28134 6976
rect 28092 6866 28120 6967
rect 27804 6860 27856 6866
rect 27804 6802 27856 6808
rect 27988 6860 28040 6866
rect 27988 6802 28040 6808
rect 28080 6860 28132 6866
rect 28080 6802 28132 6808
rect 27528 6724 27580 6730
rect 27528 6666 27580 6672
rect 27158 5879 27160 5888
rect 27212 5879 27214 5888
rect 27252 5908 27304 5914
rect 27160 5850 27212 5856
rect 27252 5850 27304 5856
rect 27540 5794 27568 6666
rect 27816 6390 27844 6802
rect 27804 6384 27856 6390
rect 27804 6326 27856 6332
rect 27264 5778 27568 5794
rect 26976 5772 27028 5778
rect 26976 5714 27028 5720
rect 27252 5772 27580 5778
rect 27304 5766 27528 5772
rect 27252 5714 27304 5720
rect 27528 5714 27580 5720
rect 27712 5772 27764 5778
rect 27712 5714 27764 5720
rect 27724 5642 27752 5714
rect 27712 5636 27764 5642
rect 27712 5578 27764 5584
rect 26884 5296 26936 5302
rect 26884 5238 26936 5244
rect 26976 5296 27028 5302
rect 26976 5238 27028 5244
rect 26608 5160 26660 5166
rect 26608 5102 26660 5108
rect 26988 4758 27016 5238
rect 27712 5092 27764 5098
rect 27712 5034 27764 5040
rect 26976 4752 27028 4758
rect 26976 4694 27028 4700
rect 25464 4644 25544 4672
rect 26424 4684 26476 4690
rect 25412 4626 25464 4632
rect 26424 4626 26476 4632
rect 26056 4072 26108 4078
rect 26056 4014 26108 4020
rect 25504 3732 25556 3738
rect 25504 3674 25556 3680
rect 24952 2304 25004 2310
rect 24952 2246 25004 2252
rect 25516 800 25544 3674
rect 26068 3194 26096 4014
rect 26804 4010 26924 4026
rect 26792 4004 26924 4010
rect 26844 3998 26924 4004
rect 26792 3946 26844 3952
rect 26790 3904 26846 3913
rect 26790 3839 26846 3848
rect 26240 3528 26292 3534
rect 26240 3470 26292 3476
rect 26056 3188 26108 3194
rect 26056 3130 26108 3136
rect 26068 2582 26096 3130
rect 26252 2922 26280 3470
rect 26804 3369 26832 3839
rect 26790 3360 26846 3369
rect 26790 3295 26846 3304
rect 26330 2952 26386 2961
rect 26240 2916 26292 2922
rect 26330 2887 26386 2896
rect 26240 2858 26292 2864
rect 26056 2576 26108 2582
rect 26056 2518 26108 2524
rect 26344 800 26372 2887
rect 26896 2514 26924 3998
rect 27252 3936 27304 3942
rect 27252 3878 27304 3884
rect 27344 3936 27396 3942
rect 27344 3878 27396 3884
rect 26974 3632 27030 3641
rect 26974 3567 27030 3576
rect 26988 2825 27016 3567
rect 26974 2816 27030 2825
rect 26974 2751 27030 2760
rect 26884 2508 26936 2514
rect 26884 2450 26936 2456
rect 27264 1578 27292 3878
rect 27356 3738 27384 3878
rect 27344 3732 27396 3738
rect 27344 3674 27396 3680
rect 27724 3670 27752 5034
rect 27816 4282 27844 6326
rect 28000 5846 28028 6802
rect 27988 5840 28040 5846
rect 27988 5782 28040 5788
rect 28184 4826 28212 15030
rect 28816 14816 28868 14822
rect 28816 14758 28868 14764
rect 28264 13320 28316 13326
rect 28264 13262 28316 13268
rect 28448 13320 28500 13326
rect 28448 13262 28500 13268
rect 28276 12170 28304 13262
rect 28460 12850 28488 13262
rect 28724 13184 28776 13190
rect 28724 13126 28776 13132
rect 28448 12844 28500 12850
rect 28448 12786 28500 12792
rect 28540 12776 28592 12782
rect 28540 12718 28592 12724
rect 28264 12164 28316 12170
rect 28264 12106 28316 12112
rect 28356 11824 28408 11830
rect 28356 11766 28408 11772
rect 28264 11280 28316 11286
rect 28264 11222 28316 11228
rect 28276 6866 28304 11222
rect 28368 11218 28396 11766
rect 28356 11212 28408 11218
rect 28552 11200 28580 12718
rect 28736 12306 28764 13126
rect 28828 12306 28856 14758
rect 28920 14550 28948 15524
rect 28908 14544 28960 14550
rect 28908 14486 28960 14492
rect 28908 14340 28960 14346
rect 28908 14282 28960 14288
rect 28724 12300 28776 12306
rect 28724 12242 28776 12248
rect 28816 12300 28868 12306
rect 28816 12242 28868 12248
rect 28356 11154 28408 11160
rect 28460 11172 28580 11200
rect 28264 6860 28316 6866
rect 28264 6802 28316 6808
rect 28264 6452 28316 6458
rect 28264 6394 28316 6400
rect 28276 5545 28304 6394
rect 28356 6384 28408 6390
rect 28356 6326 28408 6332
rect 28368 5846 28396 6326
rect 28356 5840 28408 5846
rect 28356 5782 28408 5788
rect 28262 5536 28318 5545
rect 28262 5471 28318 5480
rect 28460 5302 28488 11172
rect 28630 10568 28686 10577
rect 28630 10503 28686 10512
rect 28540 6860 28592 6866
rect 28540 6802 28592 6808
rect 28552 6497 28580 6802
rect 28538 6488 28594 6497
rect 28538 6423 28594 6432
rect 28448 5296 28500 5302
rect 28448 5238 28500 5244
rect 28172 4820 28224 4826
rect 28172 4762 28224 4768
rect 28644 4622 28672 10503
rect 28920 9110 28948 14282
rect 29288 14074 29316 15982
rect 29564 15638 29592 15982
rect 29552 15632 29604 15638
rect 29552 15574 29604 15580
rect 32876 15502 32904 16526
rect 33876 16040 33928 16046
rect 33876 15982 33928 15988
rect 33888 15706 33916 15982
rect 33876 15700 33928 15706
rect 33876 15642 33928 15648
rect 32864 15496 32916 15502
rect 32864 15438 32916 15444
rect 33140 15496 33192 15502
rect 33140 15438 33192 15444
rect 31116 15360 31168 15366
rect 31116 15302 31168 15308
rect 33048 15360 33100 15366
rect 33048 15302 33100 15308
rect 30932 14952 30984 14958
rect 30932 14894 30984 14900
rect 30748 14884 30800 14890
rect 30748 14826 30800 14832
rect 30656 14816 30708 14822
rect 30656 14758 30708 14764
rect 29460 14476 29512 14482
rect 29460 14418 29512 14424
rect 29472 14074 29500 14418
rect 29276 14068 29328 14074
rect 29276 14010 29328 14016
rect 29460 14068 29512 14074
rect 29460 14010 29512 14016
rect 29288 13938 29316 14010
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 30472 13864 30524 13870
rect 30472 13806 30524 13812
rect 30288 13796 30340 13802
rect 30288 13738 30340 13744
rect 30104 13252 30156 13258
rect 30104 13194 30156 13200
rect 29366 12744 29422 12753
rect 29366 12679 29368 12688
rect 29420 12679 29422 12688
rect 29368 12650 29420 12656
rect 29644 12640 29696 12646
rect 29644 12582 29696 12588
rect 29656 12374 29684 12582
rect 30010 12472 30066 12481
rect 30010 12407 30012 12416
rect 30064 12407 30066 12416
rect 30012 12378 30064 12384
rect 30116 12374 30144 13194
rect 30300 13190 30328 13738
rect 30380 13388 30432 13394
rect 30380 13330 30432 13336
rect 30288 13184 30340 13190
rect 30288 13126 30340 13132
rect 29644 12368 29696 12374
rect 29644 12310 29696 12316
rect 30104 12368 30156 12374
rect 30104 12310 30156 12316
rect 29828 11620 29880 11626
rect 29828 11562 29880 11568
rect 29840 11354 29868 11562
rect 29828 11348 29880 11354
rect 29828 11290 29880 11296
rect 29000 11212 29052 11218
rect 29000 11154 29052 11160
rect 29012 11082 29040 11154
rect 29000 11076 29052 11082
rect 29000 11018 29052 11024
rect 29012 10130 29040 11018
rect 30116 10606 30144 12310
rect 30196 12300 30248 12306
rect 30196 12242 30248 12248
rect 30208 11830 30236 12242
rect 30196 11824 30248 11830
rect 30196 11766 30248 11772
rect 30196 11688 30248 11694
rect 30196 11630 30248 11636
rect 30208 11218 30236 11630
rect 30196 11212 30248 11218
rect 30196 11154 30248 11160
rect 30104 10600 30156 10606
rect 30104 10542 30156 10548
rect 29736 10260 29788 10266
rect 29736 10202 29788 10208
rect 29000 10124 29052 10130
rect 29000 10066 29052 10072
rect 29012 9518 29040 10066
rect 29748 9586 29776 10202
rect 29736 9580 29788 9586
rect 29736 9522 29788 9528
rect 29000 9512 29052 9518
rect 29000 9454 29052 9460
rect 29276 9444 29328 9450
rect 29276 9386 29328 9392
rect 28908 9104 28960 9110
rect 28908 9046 28960 9052
rect 29184 9036 29236 9042
rect 29184 8978 29236 8984
rect 29000 7948 29052 7954
rect 29000 7890 29052 7896
rect 29012 7342 29040 7890
rect 29000 7336 29052 7342
rect 29000 7278 29052 7284
rect 29012 7206 29040 7278
rect 29000 7200 29052 7206
rect 29000 7142 29052 7148
rect 28724 6792 28776 6798
rect 28724 6734 28776 6740
rect 28736 5030 28764 6734
rect 29196 6338 29224 8978
rect 28920 6310 29224 6338
rect 28920 6254 28948 6310
rect 28908 6248 28960 6254
rect 28908 6190 28960 6196
rect 28816 5568 28868 5574
rect 28814 5536 28816 5545
rect 29092 5568 29144 5574
rect 28868 5536 28870 5545
rect 29092 5510 29144 5516
rect 28814 5471 28870 5480
rect 28724 5024 28776 5030
rect 28724 4966 28776 4972
rect 28632 4616 28684 4622
rect 28632 4558 28684 4564
rect 28736 4486 28764 4966
rect 29000 4820 29052 4826
rect 29000 4762 29052 4768
rect 28908 4548 28960 4554
rect 28908 4490 28960 4496
rect 28356 4480 28408 4486
rect 28356 4422 28408 4428
rect 28724 4480 28776 4486
rect 28724 4422 28776 4428
rect 27804 4276 27856 4282
rect 27804 4218 27856 4224
rect 27816 3738 27844 4218
rect 28264 4140 28316 4146
rect 28264 4082 28316 4088
rect 27804 3732 27856 3738
rect 27804 3674 27856 3680
rect 28276 3670 28304 4082
rect 27712 3664 27764 3670
rect 27342 3632 27398 3641
rect 27712 3606 27764 3612
rect 27896 3664 27948 3670
rect 27896 3606 27948 3612
rect 28264 3664 28316 3670
rect 28264 3606 28316 3612
rect 27342 3567 27398 3576
rect 27172 1550 27292 1578
rect 27172 1358 27200 1550
rect 27356 1442 27384 3567
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 27540 3126 27568 3470
rect 27528 3120 27580 3126
rect 27528 3062 27580 3068
rect 27908 2990 27936 3606
rect 28080 3188 28132 3194
rect 28080 3130 28132 3136
rect 27896 2984 27948 2990
rect 27896 2926 27948 2932
rect 27264 1414 27384 1442
rect 27160 1352 27212 1358
rect 27160 1294 27212 1300
rect 27264 800 27292 1414
rect 28092 800 28120 3130
rect 28276 2514 28304 3606
rect 28368 3058 28396 4422
rect 28920 4282 28948 4490
rect 28908 4276 28960 4282
rect 28908 4218 28960 4224
rect 29012 4078 29040 4762
rect 29104 4758 29132 5510
rect 29092 4752 29144 4758
rect 29092 4694 29144 4700
rect 29196 4690 29224 6310
rect 29288 6118 29316 9386
rect 29736 8832 29788 8838
rect 29736 8774 29788 8780
rect 30196 8832 30248 8838
rect 30196 8774 30248 8780
rect 29748 8430 29776 8774
rect 29552 8424 29604 8430
rect 29552 8366 29604 8372
rect 29736 8424 29788 8430
rect 29736 8366 29788 8372
rect 29564 7342 29592 8366
rect 29552 7336 29604 7342
rect 29552 7278 29604 7284
rect 29460 6656 29512 6662
rect 29460 6598 29512 6604
rect 29472 6254 29500 6598
rect 29368 6248 29420 6254
rect 29368 6190 29420 6196
rect 29460 6248 29512 6254
rect 29460 6190 29512 6196
rect 29276 6112 29328 6118
rect 29276 6054 29328 6060
rect 29288 5710 29316 6054
rect 29276 5704 29328 5710
rect 29276 5646 29328 5652
rect 29380 5545 29408 6190
rect 29472 6118 29500 6190
rect 29460 6112 29512 6118
rect 29460 6054 29512 6060
rect 29366 5536 29422 5545
rect 29366 5471 29422 5480
rect 29184 4684 29236 4690
rect 29184 4626 29236 4632
rect 29000 4072 29052 4078
rect 29000 4014 29052 4020
rect 29276 4072 29328 4078
rect 29276 4014 29328 4020
rect 29288 3398 29316 4014
rect 29380 3398 29408 5471
rect 29564 4078 29592 7278
rect 30208 7177 30236 8774
rect 30392 8498 30420 13330
rect 30484 13258 30512 13806
rect 30472 13252 30524 13258
rect 30472 13194 30524 13200
rect 30668 12782 30696 14758
rect 30760 13870 30788 14826
rect 30840 14476 30892 14482
rect 30840 14418 30892 14424
rect 30748 13864 30800 13870
rect 30748 13806 30800 13812
rect 30760 13394 30788 13806
rect 30748 13388 30800 13394
rect 30748 13330 30800 13336
rect 30852 12986 30880 14418
rect 30944 14278 30972 14894
rect 31128 14550 31156 15302
rect 31500 15260 31796 15280
rect 31556 15258 31580 15260
rect 31636 15258 31660 15260
rect 31716 15258 31740 15260
rect 31578 15206 31580 15258
rect 31642 15206 31654 15258
rect 31716 15206 31718 15258
rect 31556 15204 31580 15206
rect 31636 15204 31660 15206
rect 31716 15204 31740 15206
rect 31500 15184 31796 15204
rect 33060 15162 33088 15302
rect 33152 15162 33180 15438
rect 33888 15434 33916 15642
rect 33876 15428 33928 15434
rect 33876 15370 33928 15376
rect 33048 15156 33100 15162
rect 33048 15098 33100 15104
rect 33140 15156 33192 15162
rect 33140 15098 33192 15104
rect 32864 14952 32916 14958
rect 32864 14894 32916 14900
rect 31116 14544 31168 14550
rect 31116 14486 31168 14492
rect 30932 14272 30984 14278
rect 30932 14214 30984 14220
rect 32496 14272 32548 14278
rect 32496 14214 32548 14220
rect 31500 14172 31796 14192
rect 31556 14170 31580 14172
rect 31636 14170 31660 14172
rect 31716 14170 31740 14172
rect 31578 14118 31580 14170
rect 31642 14118 31654 14170
rect 31716 14118 31718 14170
rect 31556 14116 31580 14118
rect 31636 14116 31660 14118
rect 31716 14116 31740 14118
rect 31500 14096 31796 14116
rect 31116 13728 31168 13734
rect 31116 13670 31168 13676
rect 31128 13258 31156 13670
rect 32036 13456 32088 13462
rect 32036 13398 32088 13404
rect 31116 13252 31168 13258
rect 31116 13194 31168 13200
rect 30932 13184 30984 13190
rect 30932 13126 30984 13132
rect 30840 12980 30892 12986
rect 30840 12922 30892 12928
rect 30656 12776 30708 12782
rect 30656 12718 30708 12724
rect 30748 12368 30800 12374
rect 30748 12310 30800 12316
rect 30472 12232 30524 12238
rect 30470 12200 30472 12209
rect 30524 12200 30526 12209
rect 30470 12135 30526 12144
rect 30760 11762 30788 12310
rect 30748 11756 30800 11762
rect 30748 11698 30800 11704
rect 30668 11626 30880 11642
rect 30656 11620 30880 11626
rect 30708 11614 30880 11620
rect 30656 11562 30708 11568
rect 30852 11558 30880 11614
rect 30840 11552 30892 11558
rect 30840 11494 30892 11500
rect 30944 11354 30972 13126
rect 31500 13084 31796 13104
rect 31556 13082 31580 13084
rect 31636 13082 31660 13084
rect 31716 13082 31740 13084
rect 31578 13030 31580 13082
rect 31642 13030 31654 13082
rect 31716 13030 31718 13082
rect 31556 13028 31580 13030
rect 31636 13028 31660 13030
rect 31716 13028 31740 13030
rect 31500 13008 31796 13028
rect 32048 12986 32076 13398
rect 32404 13388 32456 13394
rect 32404 13330 32456 13336
rect 32036 12980 32088 12986
rect 32036 12922 32088 12928
rect 32416 12374 32444 13330
rect 31024 12368 31076 12374
rect 31024 12310 31076 12316
rect 32404 12368 32456 12374
rect 32404 12310 32456 12316
rect 31036 12170 31064 12310
rect 32220 12300 32272 12306
rect 32220 12242 32272 12248
rect 31208 12232 31260 12238
rect 31206 12200 31208 12209
rect 31260 12200 31262 12209
rect 31024 12164 31076 12170
rect 31206 12135 31262 12144
rect 31024 12106 31076 12112
rect 31500 11996 31796 12016
rect 31556 11994 31580 11996
rect 31636 11994 31660 11996
rect 31716 11994 31740 11996
rect 31578 11942 31580 11994
rect 31642 11942 31654 11994
rect 31716 11942 31718 11994
rect 31556 11940 31580 11942
rect 31636 11940 31660 11942
rect 31716 11940 31740 11942
rect 31500 11920 31796 11940
rect 32232 11694 32260 12242
rect 32404 11892 32456 11898
rect 32404 11834 32456 11840
rect 32416 11694 32444 11834
rect 32508 11744 32536 14214
rect 32876 13870 32904 14894
rect 33060 14550 33088 15098
rect 33324 14952 33376 14958
rect 33324 14894 33376 14900
rect 33048 14544 33100 14550
rect 33048 14486 33100 14492
rect 33336 14074 33364 14894
rect 33416 14884 33468 14890
rect 33416 14826 33468 14832
rect 33428 14550 33456 14826
rect 34256 14550 34284 16934
rect 34796 16652 34848 16658
rect 34796 16594 34848 16600
rect 34612 14816 34664 14822
rect 34612 14758 34664 14764
rect 33416 14544 33468 14550
rect 33416 14486 33468 14492
rect 34244 14544 34296 14550
rect 34244 14486 34296 14492
rect 34624 14482 34652 14758
rect 34612 14476 34664 14482
rect 34612 14418 34664 14424
rect 34808 14278 34836 16594
rect 34900 16250 34928 16934
rect 35452 16810 35480 18835
rect 37384 17218 37412 18835
rect 37292 17202 37412 17218
rect 37280 17196 37412 17202
rect 37332 17190 37412 17196
rect 37280 17138 37332 17144
rect 35992 17060 36044 17066
rect 35992 17002 36044 17008
rect 36820 17060 36872 17066
rect 36820 17002 36872 17008
rect 35452 16782 35572 16810
rect 35164 16652 35216 16658
rect 35164 16594 35216 16600
rect 34888 16244 34940 16250
rect 34888 16186 34940 16192
rect 34900 16046 34928 16186
rect 34888 16040 34940 16046
rect 34888 15982 34940 15988
rect 35176 15162 35204 16594
rect 35544 16590 35572 16782
rect 35256 16584 35308 16590
rect 35256 16526 35308 16532
rect 35532 16584 35584 16590
rect 35532 16526 35584 16532
rect 35268 16114 35296 16526
rect 35256 16108 35308 16114
rect 35256 16050 35308 16056
rect 35544 16046 35572 16526
rect 35532 16040 35584 16046
rect 35532 15982 35584 15988
rect 35348 15972 35400 15978
rect 35348 15914 35400 15920
rect 35164 15156 35216 15162
rect 35164 15098 35216 15104
rect 35360 14958 35388 15914
rect 36004 15638 36032 17002
rect 36832 16794 36860 17002
rect 36820 16788 36872 16794
rect 36820 16730 36872 16736
rect 37384 16250 37412 17190
rect 38936 17196 38988 17202
rect 38936 17138 38988 17144
rect 37832 17128 37884 17134
rect 37832 17070 37884 17076
rect 38752 17128 38804 17134
rect 38752 17070 38804 17076
rect 37844 16658 37872 17070
rect 37832 16652 37884 16658
rect 37832 16594 37884 16600
rect 37372 16244 37424 16250
rect 37372 16186 37424 16192
rect 37844 16114 37872 16594
rect 37832 16108 37884 16114
rect 37832 16050 37884 16056
rect 36544 16040 36596 16046
rect 36544 15982 36596 15988
rect 36084 15700 36136 15706
rect 36084 15642 36136 15648
rect 35992 15632 36044 15638
rect 35992 15574 36044 15580
rect 36096 15502 36124 15642
rect 36176 15564 36228 15570
rect 36176 15506 36228 15512
rect 36084 15496 36136 15502
rect 36084 15438 36136 15444
rect 36096 15026 36124 15438
rect 36188 15094 36216 15506
rect 36556 15366 36584 15982
rect 37740 15564 37792 15570
rect 37740 15506 37792 15512
rect 36544 15360 36596 15366
rect 36544 15302 36596 15308
rect 37372 15156 37424 15162
rect 37372 15098 37424 15104
rect 36176 15088 36228 15094
rect 36176 15030 36228 15036
rect 37384 15026 37412 15098
rect 36084 15020 36136 15026
rect 36084 14962 36136 14968
rect 37372 15020 37424 15026
rect 37372 14962 37424 14968
rect 35348 14952 35400 14958
rect 35348 14894 35400 14900
rect 35716 14476 35768 14482
rect 35716 14418 35768 14424
rect 34796 14272 34848 14278
rect 34796 14214 34848 14220
rect 34888 14272 34940 14278
rect 34888 14214 34940 14220
rect 33324 14068 33376 14074
rect 33324 14010 33376 14016
rect 32864 13864 32916 13870
rect 32864 13806 32916 13812
rect 34900 13462 34928 14214
rect 35164 13796 35216 13802
rect 35164 13738 35216 13744
rect 34888 13456 34940 13462
rect 34888 13398 34940 13404
rect 35176 13394 35204 13738
rect 35164 13388 35216 13394
rect 35164 13330 35216 13336
rect 33876 13320 33928 13326
rect 33876 13262 33928 13268
rect 35072 13320 35124 13326
rect 35072 13262 35124 13268
rect 33692 13184 33744 13190
rect 33692 13126 33744 13132
rect 33784 13184 33836 13190
rect 33784 13126 33836 13132
rect 32588 12776 32640 12782
rect 32588 12718 32640 12724
rect 32956 12776 33008 12782
rect 32956 12718 33008 12724
rect 32600 12238 32628 12718
rect 32968 12374 32996 12718
rect 33508 12708 33560 12714
rect 33508 12650 33560 12656
rect 32956 12368 33008 12374
rect 32956 12310 33008 12316
rect 32772 12300 32824 12306
rect 32772 12242 32824 12248
rect 32588 12232 32640 12238
rect 32588 12174 32640 12180
rect 32588 11756 32640 11762
rect 32508 11716 32588 11744
rect 32588 11698 32640 11704
rect 32220 11688 32272 11694
rect 32220 11630 32272 11636
rect 32404 11688 32456 11694
rect 32404 11630 32456 11636
rect 32784 11626 32812 12242
rect 33520 11694 33548 12650
rect 33704 11762 33732 13126
rect 33796 12238 33824 13126
rect 33888 12889 33916 13262
rect 34244 13184 34296 13190
rect 34244 13126 34296 13132
rect 33874 12880 33930 12889
rect 33874 12815 33930 12824
rect 33784 12232 33836 12238
rect 33784 12174 33836 12180
rect 33692 11756 33744 11762
rect 33888 11744 33916 12815
rect 34256 12753 34284 13126
rect 34428 12844 34480 12850
rect 34428 12786 34480 12792
rect 34242 12744 34298 12753
rect 34242 12679 34298 12688
rect 34336 12300 34388 12306
rect 34336 12242 34388 12248
rect 33968 12232 34020 12238
rect 33968 12174 34020 12180
rect 33980 11762 34008 12174
rect 34244 12096 34296 12102
rect 34244 12038 34296 12044
rect 33692 11698 33744 11704
rect 33796 11716 33916 11744
rect 33968 11756 34020 11762
rect 33508 11688 33560 11694
rect 33508 11630 33560 11636
rect 32772 11620 32824 11626
rect 32772 11562 32824 11568
rect 30932 11348 30984 11354
rect 30932 11290 30984 11296
rect 31116 11348 31168 11354
rect 31116 11290 31168 11296
rect 32312 11348 32364 11354
rect 32312 11290 32364 11296
rect 30472 11212 30524 11218
rect 30472 11154 30524 11160
rect 30484 10538 30512 11154
rect 30656 10600 30708 10606
rect 30656 10542 30708 10548
rect 30472 10532 30524 10538
rect 30472 10474 30524 10480
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 30484 7206 30512 10474
rect 30668 10130 30696 10542
rect 30840 10464 30892 10470
rect 30840 10406 30892 10412
rect 30656 10124 30708 10130
rect 30656 10066 30708 10072
rect 30748 9444 30800 9450
rect 30748 9386 30800 9392
rect 30760 9178 30788 9386
rect 30748 9172 30800 9178
rect 30748 9114 30800 9120
rect 30656 9036 30708 9042
rect 30656 8978 30708 8984
rect 30564 8832 30616 8838
rect 30564 8774 30616 8780
rect 30472 7200 30524 7206
rect 30194 7168 30250 7177
rect 30472 7142 30524 7148
rect 30194 7103 30250 7112
rect 30012 6656 30064 6662
rect 30012 6598 30064 6604
rect 30104 6656 30156 6662
rect 30104 6598 30156 6604
rect 30024 6118 30052 6598
rect 30012 6112 30064 6118
rect 30012 6054 30064 6060
rect 30116 5778 30144 6598
rect 30208 5846 30236 7103
rect 30576 6866 30604 8774
rect 30668 8294 30696 8978
rect 30852 8566 30880 10406
rect 30840 8560 30892 8566
rect 30840 8502 30892 8508
rect 31024 8424 31076 8430
rect 31024 8366 31076 8372
rect 30656 8288 30708 8294
rect 30656 8230 30708 8236
rect 30668 6866 30696 8230
rect 30840 7200 30892 7206
rect 30840 7142 30892 7148
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30656 6860 30708 6866
rect 30656 6802 30708 6808
rect 30472 6180 30524 6186
rect 30472 6122 30524 6128
rect 30286 6080 30342 6089
rect 30286 6015 30342 6024
rect 30196 5840 30248 5846
rect 30196 5782 30248 5788
rect 30104 5772 30156 5778
rect 30104 5714 30156 5720
rect 30196 5704 30248 5710
rect 30196 5646 30248 5652
rect 30208 4865 30236 5646
rect 30194 4856 30250 4865
rect 30194 4791 30250 4800
rect 29736 4684 29788 4690
rect 29736 4626 29788 4632
rect 29552 4072 29604 4078
rect 29552 4014 29604 4020
rect 29748 3670 29776 4626
rect 30104 4004 30156 4010
rect 30104 3946 30156 3952
rect 30116 3738 30144 3946
rect 30104 3732 30156 3738
rect 30104 3674 30156 3680
rect 29736 3664 29788 3670
rect 29736 3606 29788 3612
rect 29276 3392 29328 3398
rect 29276 3334 29328 3340
rect 29368 3392 29420 3398
rect 29368 3334 29420 3340
rect 28356 3052 28408 3058
rect 28356 2994 28408 3000
rect 29000 3052 29052 3058
rect 29000 2994 29052 3000
rect 28264 2508 28316 2514
rect 28264 2450 28316 2456
rect 29012 800 29040 2994
rect 29748 2310 29776 3606
rect 30012 3596 30064 3602
rect 30012 3538 30064 3544
rect 29826 3088 29882 3097
rect 29826 3023 29882 3032
rect 29736 2304 29788 2310
rect 29736 2246 29788 2252
rect 29840 800 29868 3023
rect 30024 2990 30052 3538
rect 30300 3058 30328 6015
rect 30484 5710 30512 6122
rect 30472 5704 30524 5710
rect 30576 5681 30604 6802
rect 30472 5646 30524 5652
rect 30562 5672 30618 5681
rect 30484 3058 30512 5646
rect 30562 5607 30618 5616
rect 30564 5024 30616 5030
rect 30564 4966 30616 4972
rect 30576 4622 30604 4966
rect 30852 4826 30880 7142
rect 30932 6180 30984 6186
rect 30932 6122 30984 6128
rect 30944 5914 30972 6122
rect 30932 5908 30984 5914
rect 30932 5850 30984 5856
rect 30930 5808 30986 5817
rect 30930 5743 30932 5752
rect 30984 5743 30986 5752
rect 30932 5714 30984 5720
rect 30840 4820 30892 4826
rect 30840 4762 30892 4768
rect 31036 4690 31064 8366
rect 31128 5778 31156 11290
rect 31500 10908 31796 10928
rect 31556 10906 31580 10908
rect 31636 10906 31660 10908
rect 31716 10906 31740 10908
rect 31578 10854 31580 10906
rect 31642 10854 31654 10906
rect 31716 10854 31718 10906
rect 31556 10852 31580 10854
rect 31636 10852 31660 10854
rect 31716 10852 31740 10854
rect 31500 10832 31796 10852
rect 32324 10810 32352 11290
rect 33508 11144 33560 11150
rect 33508 11086 33560 11092
rect 32312 10804 32364 10810
rect 32312 10746 32364 10752
rect 31852 10600 31904 10606
rect 31852 10542 31904 10548
rect 33140 10600 33192 10606
rect 33140 10542 33192 10548
rect 31500 9820 31796 9840
rect 31556 9818 31580 9820
rect 31636 9818 31660 9820
rect 31716 9818 31740 9820
rect 31578 9766 31580 9818
rect 31642 9766 31654 9818
rect 31716 9766 31718 9818
rect 31556 9764 31580 9766
rect 31636 9764 31660 9766
rect 31716 9764 31740 9766
rect 31298 9752 31354 9761
rect 31500 9744 31796 9764
rect 31298 9687 31354 9696
rect 31312 9382 31340 9687
rect 31864 9518 31892 10542
rect 32036 10464 32088 10470
rect 32036 10406 32088 10412
rect 31852 9512 31904 9518
rect 31852 9454 31904 9460
rect 31300 9376 31352 9382
rect 31300 9318 31352 9324
rect 31300 8968 31352 8974
rect 31300 8910 31352 8916
rect 31312 6254 31340 8910
rect 31500 8732 31796 8752
rect 31556 8730 31580 8732
rect 31636 8730 31660 8732
rect 31716 8730 31740 8732
rect 31578 8678 31580 8730
rect 31642 8678 31654 8730
rect 31716 8678 31718 8730
rect 31556 8676 31580 8678
rect 31636 8676 31660 8678
rect 31716 8676 31740 8678
rect 31500 8656 31796 8676
rect 32048 8634 32076 10406
rect 32128 10124 32180 10130
rect 32128 10066 32180 10072
rect 32312 10124 32364 10130
rect 32312 10066 32364 10072
rect 32140 9042 32168 10066
rect 32220 10056 32272 10062
rect 32220 9998 32272 10004
rect 32128 9036 32180 9042
rect 32128 8978 32180 8984
rect 32036 8628 32088 8634
rect 32036 8570 32088 8576
rect 31850 8528 31906 8537
rect 31850 8463 31852 8472
rect 31904 8463 31906 8472
rect 32126 8528 32182 8537
rect 32126 8463 32182 8472
rect 31852 8434 31904 8440
rect 31944 8016 31996 8022
rect 31944 7958 31996 7964
rect 31392 7880 31444 7886
rect 31392 7822 31444 7828
rect 31404 7478 31432 7822
rect 31500 7644 31796 7664
rect 31556 7642 31580 7644
rect 31636 7642 31660 7644
rect 31716 7642 31740 7644
rect 31578 7590 31580 7642
rect 31642 7590 31654 7642
rect 31716 7590 31718 7642
rect 31556 7588 31580 7590
rect 31636 7588 31660 7590
rect 31716 7588 31740 7590
rect 31500 7568 31796 7588
rect 31956 7478 31984 7958
rect 32036 7948 32088 7954
rect 32036 7890 32088 7896
rect 31392 7472 31444 7478
rect 31392 7414 31444 7420
rect 31944 7472 31996 7478
rect 31944 7414 31996 7420
rect 31208 6248 31260 6254
rect 31206 6216 31208 6225
rect 31300 6248 31352 6254
rect 31260 6216 31262 6225
rect 31300 6190 31352 6196
rect 31206 6151 31262 6160
rect 31312 6100 31340 6190
rect 31220 6072 31340 6100
rect 31116 5772 31168 5778
rect 31116 5714 31168 5720
rect 31116 4752 31168 4758
rect 31116 4694 31168 4700
rect 31024 4684 31076 4690
rect 31024 4626 31076 4632
rect 30564 4616 30616 4622
rect 30564 4558 30616 4564
rect 31022 4584 31078 4593
rect 30576 3466 30604 4558
rect 31022 4519 31078 4528
rect 31036 4486 31064 4519
rect 31024 4480 31076 4486
rect 31024 4422 31076 4428
rect 31024 4072 31076 4078
rect 30654 4040 30710 4049
rect 31024 4014 31076 4020
rect 30654 3975 30710 3984
rect 30932 4004 30984 4010
rect 30564 3460 30616 3466
rect 30564 3402 30616 3408
rect 30288 3052 30340 3058
rect 30288 2994 30340 3000
rect 30472 3052 30524 3058
rect 30472 2994 30524 3000
rect 30012 2984 30064 2990
rect 30012 2926 30064 2932
rect 30024 2650 30052 2926
rect 30288 2916 30340 2922
rect 30288 2858 30340 2864
rect 30380 2916 30432 2922
rect 30380 2858 30432 2864
rect 30012 2644 30064 2650
rect 30012 2586 30064 2592
rect 30300 2514 30328 2858
rect 30392 2689 30420 2858
rect 30378 2680 30434 2689
rect 30378 2615 30434 2624
rect 30288 2508 30340 2514
rect 30288 2450 30340 2456
rect 30668 800 30696 3975
rect 30932 3946 30984 3952
rect 30748 3460 30800 3466
rect 30748 3402 30800 3408
rect 30760 2990 30788 3402
rect 30944 3058 30972 3946
rect 31036 3058 31064 4014
rect 31128 4010 31156 4694
rect 31220 4146 31248 6072
rect 31298 5944 31354 5953
rect 31298 5879 31300 5888
rect 31352 5879 31354 5888
rect 31300 5850 31352 5856
rect 31300 4480 31352 4486
rect 31300 4422 31352 4428
rect 31208 4140 31260 4146
rect 31208 4082 31260 4088
rect 31312 4078 31340 4422
rect 31404 4282 31432 7414
rect 32048 7041 32076 7890
rect 32034 7032 32090 7041
rect 32140 7018 32168 8463
rect 32232 7993 32260 9998
rect 32324 9178 32352 10066
rect 32404 9580 32456 9586
rect 32404 9522 32456 9528
rect 32416 9382 32444 9522
rect 32680 9512 32732 9518
rect 32680 9454 32732 9460
rect 32404 9376 32456 9382
rect 32404 9318 32456 9324
rect 32312 9172 32364 9178
rect 32312 9114 32364 9120
rect 32324 8430 32352 9114
rect 32496 9036 32548 9042
rect 32496 8978 32548 8984
rect 32312 8424 32364 8430
rect 32312 8366 32364 8372
rect 32218 7984 32274 7993
rect 32218 7919 32274 7928
rect 32324 7750 32352 8366
rect 32404 7880 32456 7886
rect 32404 7822 32456 7828
rect 32312 7744 32364 7750
rect 32312 7686 32364 7692
rect 32140 6990 32260 7018
rect 32034 6967 32090 6976
rect 32048 6916 32076 6967
rect 32048 6888 32168 6916
rect 31500 6556 31796 6576
rect 31556 6554 31580 6556
rect 31636 6554 31660 6556
rect 31716 6554 31740 6556
rect 31578 6502 31580 6554
rect 31642 6502 31654 6554
rect 31716 6502 31718 6554
rect 31556 6500 31580 6502
rect 31636 6500 31660 6502
rect 31716 6500 31740 6502
rect 31500 6480 31796 6500
rect 31760 6248 31812 6254
rect 31760 6190 31812 6196
rect 31772 6089 31800 6190
rect 31758 6080 31814 6089
rect 31758 6015 31814 6024
rect 31850 5672 31906 5681
rect 31850 5607 31852 5616
rect 31904 5607 31906 5616
rect 31852 5578 31904 5584
rect 31500 5468 31796 5488
rect 31556 5466 31580 5468
rect 31636 5466 31660 5468
rect 31716 5466 31740 5468
rect 31578 5414 31580 5466
rect 31642 5414 31654 5466
rect 31716 5414 31718 5466
rect 31556 5412 31580 5414
rect 31636 5412 31660 5414
rect 31716 5412 31740 5414
rect 31500 5392 31796 5412
rect 31944 5160 31996 5166
rect 31944 5102 31996 5108
rect 31956 4826 31984 5102
rect 31944 4820 31996 4826
rect 31944 4762 31996 4768
rect 31944 4684 31996 4690
rect 31944 4626 31996 4632
rect 32036 4684 32088 4690
rect 32036 4626 32088 4632
rect 31500 4380 31796 4400
rect 31556 4378 31580 4380
rect 31636 4378 31660 4380
rect 31716 4378 31740 4380
rect 31578 4326 31580 4378
rect 31642 4326 31654 4378
rect 31716 4326 31718 4378
rect 31556 4324 31580 4326
rect 31636 4324 31660 4326
rect 31716 4324 31740 4326
rect 31500 4304 31796 4324
rect 31392 4276 31444 4282
rect 31392 4218 31444 4224
rect 31300 4072 31352 4078
rect 31300 4014 31352 4020
rect 31956 4026 31984 4626
rect 32048 4486 32076 4626
rect 32036 4480 32088 4486
rect 32036 4422 32088 4428
rect 31116 4004 31168 4010
rect 31956 3998 32076 4026
rect 31116 3946 31168 3952
rect 32048 3942 32076 3998
rect 31852 3936 31904 3942
rect 31852 3878 31904 3884
rect 32036 3936 32088 3942
rect 32036 3878 32088 3884
rect 31864 3777 31892 3878
rect 31666 3768 31722 3777
rect 31666 3703 31722 3712
rect 31850 3768 31906 3777
rect 31850 3703 31906 3712
rect 31680 3618 31708 3703
rect 31680 3590 31892 3618
rect 31116 3528 31168 3534
rect 31116 3470 31168 3476
rect 30932 3052 30984 3058
rect 30932 2994 30984 3000
rect 31024 3052 31076 3058
rect 31024 2994 31076 3000
rect 30748 2984 30800 2990
rect 30748 2926 30800 2932
rect 31024 2576 31076 2582
rect 31024 2518 31076 2524
rect 31036 2106 31064 2518
rect 31128 2446 31156 3470
rect 31300 3392 31352 3398
rect 31300 3334 31352 3340
rect 31864 3346 31892 3590
rect 31942 3360 31998 3369
rect 31312 3233 31340 3334
rect 31864 3318 31942 3346
rect 31500 3292 31796 3312
rect 31942 3295 31998 3304
rect 31556 3290 31580 3292
rect 31636 3290 31660 3292
rect 31716 3290 31740 3292
rect 31578 3238 31580 3290
rect 31642 3238 31654 3290
rect 31716 3238 31718 3290
rect 31556 3236 31580 3238
rect 31636 3236 31660 3238
rect 31716 3236 31740 3238
rect 31298 3224 31354 3233
rect 31500 3216 31796 3236
rect 31298 3159 31354 3168
rect 32140 3058 32168 6888
rect 32232 5250 32260 6990
rect 32312 6860 32364 6866
rect 32312 6802 32364 6808
rect 32324 5778 32352 6802
rect 32416 6610 32444 7822
rect 32508 7546 32536 8978
rect 32588 7948 32640 7954
rect 32588 7890 32640 7896
rect 32496 7540 32548 7546
rect 32496 7482 32548 7488
rect 32508 6730 32536 7482
rect 32600 7342 32628 7890
rect 32588 7336 32640 7342
rect 32588 7278 32640 7284
rect 32496 6724 32548 6730
rect 32496 6666 32548 6672
rect 32416 6582 32536 6610
rect 32404 5840 32456 5846
rect 32402 5808 32404 5817
rect 32456 5808 32458 5817
rect 32312 5772 32364 5778
rect 32402 5743 32458 5752
rect 32312 5714 32364 5720
rect 32232 5222 32444 5250
rect 32220 5160 32272 5166
rect 32220 5102 32272 5108
rect 32312 5160 32364 5166
rect 32312 5102 32364 5108
rect 32232 4282 32260 5102
rect 32220 4276 32272 4282
rect 32220 4218 32272 4224
rect 32324 3534 32352 5102
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 32128 3052 32180 3058
rect 32128 2994 32180 3000
rect 31392 2916 31444 2922
rect 31392 2858 31444 2864
rect 31116 2440 31168 2446
rect 31116 2382 31168 2388
rect 31024 2100 31076 2106
rect 31024 2042 31076 2048
rect 31404 898 31432 2858
rect 32324 2825 32352 3470
rect 32416 3398 32444 5222
rect 32508 5166 32536 6582
rect 32600 6225 32628 7278
rect 32692 6866 32720 9454
rect 32772 9376 32824 9382
rect 32772 9318 32824 9324
rect 32784 8294 32812 9318
rect 32956 8968 33008 8974
rect 32956 8910 33008 8916
rect 32772 8288 32824 8294
rect 32772 8230 32824 8236
rect 32680 6860 32732 6866
rect 32680 6802 32732 6808
rect 32784 6769 32812 8230
rect 32968 8106 32996 8910
rect 33048 8832 33100 8838
rect 33048 8774 33100 8780
rect 33060 8634 33088 8774
rect 33048 8628 33100 8634
rect 33048 8570 33100 8576
rect 33152 8498 33180 10542
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33428 9518 33456 9998
rect 33520 9654 33548 11086
rect 33600 11008 33652 11014
rect 33600 10950 33652 10956
rect 33612 10130 33640 10950
rect 33796 10606 33824 11716
rect 33968 11698 34020 11704
rect 34152 11688 34204 11694
rect 34152 11630 34204 11636
rect 33968 11552 34020 11558
rect 33968 11494 34020 11500
rect 33980 11218 34008 11494
rect 33968 11212 34020 11218
rect 33968 11154 34020 11160
rect 33876 10736 33928 10742
rect 33876 10678 33928 10684
rect 33784 10600 33836 10606
rect 33784 10542 33836 10548
rect 33600 10124 33652 10130
rect 33600 10066 33652 10072
rect 33508 9648 33560 9654
rect 33508 9590 33560 9596
rect 33888 9518 33916 10678
rect 33416 9512 33468 9518
rect 33416 9454 33468 9460
rect 33876 9512 33928 9518
rect 33876 9454 33928 9460
rect 33416 8968 33468 8974
rect 33416 8910 33468 8916
rect 33140 8492 33192 8498
rect 33140 8434 33192 8440
rect 33232 8424 33284 8430
rect 33232 8366 33284 8372
rect 32968 8078 33180 8106
rect 32954 7984 33010 7993
rect 32954 7919 33010 7928
rect 32864 7404 32916 7410
rect 32864 7346 32916 7352
rect 32876 7313 32904 7346
rect 32862 7304 32918 7313
rect 32862 7239 32918 7248
rect 32770 6760 32826 6769
rect 32876 6730 32904 7239
rect 32770 6695 32826 6704
rect 32864 6724 32916 6730
rect 32864 6666 32916 6672
rect 32586 6216 32642 6225
rect 32586 6151 32642 6160
rect 32600 5778 32628 6151
rect 32588 5772 32640 5778
rect 32588 5714 32640 5720
rect 32680 5704 32732 5710
rect 32680 5646 32732 5652
rect 32692 5234 32720 5646
rect 32680 5228 32732 5234
rect 32680 5170 32732 5176
rect 32496 5160 32548 5166
rect 32496 5102 32548 5108
rect 32864 5092 32916 5098
rect 32864 5034 32916 5040
rect 32494 4856 32550 4865
rect 32494 4791 32550 4800
rect 32508 4690 32536 4791
rect 32496 4684 32548 4690
rect 32496 4626 32548 4632
rect 32496 4004 32548 4010
rect 32496 3946 32548 3952
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 32310 2816 32366 2825
rect 32310 2751 32366 2760
rect 31500 2204 31796 2224
rect 31556 2202 31580 2204
rect 31636 2202 31660 2204
rect 31716 2202 31740 2204
rect 31578 2150 31580 2202
rect 31642 2150 31654 2202
rect 31716 2150 31718 2202
rect 31556 2148 31580 2150
rect 31636 2148 31660 2150
rect 31716 2148 31740 2150
rect 31500 2128 31796 2148
rect 32508 898 32536 3946
rect 32680 3936 32732 3942
rect 32680 3878 32732 3884
rect 32692 2990 32720 3878
rect 32680 2984 32732 2990
rect 32680 2926 32732 2932
rect 32588 2576 32640 2582
rect 32588 2518 32640 2524
rect 32600 2106 32628 2518
rect 32772 2440 32824 2446
rect 32772 2382 32824 2388
rect 32588 2100 32640 2106
rect 32588 2042 32640 2048
rect 32784 1902 32812 2382
rect 32876 2310 32904 5034
rect 32968 4185 32996 7919
rect 33048 7268 33100 7274
rect 33048 7210 33100 7216
rect 33060 4282 33088 7210
rect 33152 4826 33180 8078
rect 33244 8022 33272 8366
rect 33428 8022 33456 8910
rect 33888 8498 33916 9454
rect 33980 9450 34008 11154
rect 34164 10130 34192 11630
rect 34256 11286 34284 12038
rect 34348 11898 34376 12242
rect 34440 12102 34468 12786
rect 34980 12232 35032 12238
rect 34980 12174 35032 12180
rect 34428 12096 34480 12102
rect 34428 12038 34480 12044
rect 34336 11892 34388 11898
rect 34336 11834 34388 11840
rect 34796 11756 34848 11762
rect 34796 11698 34848 11704
rect 34808 11626 34836 11698
rect 34796 11620 34848 11626
rect 34796 11562 34848 11568
rect 34244 11280 34296 11286
rect 34244 11222 34296 11228
rect 34992 11150 35020 12174
rect 35084 11218 35112 13262
rect 35176 12646 35204 13330
rect 35164 12640 35216 12646
rect 35164 12582 35216 12588
rect 35728 11694 35756 14418
rect 36096 14346 36124 14962
rect 36176 14952 36228 14958
rect 36176 14894 36228 14900
rect 36636 14952 36688 14958
rect 36636 14894 36688 14900
rect 36084 14340 36136 14346
rect 36084 14282 36136 14288
rect 36188 13802 36216 14894
rect 36176 13796 36228 13802
rect 36176 13738 36228 13744
rect 36176 13388 36228 13394
rect 36176 13330 36228 13336
rect 36082 12880 36138 12889
rect 36082 12815 36138 12824
rect 36096 12782 36124 12815
rect 36188 12782 36216 13330
rect 36360 13252 36412 13258
rect 36360 13194 36412 13200
rect 35900 12776 35952 12782
rect 35900 12718 35952 12724
rect 36084 12776 36136 12782
rect 36084 12718 36136 12724
rect 36176 12776 36228 12782
rect 36176 12718 36228 12724
rect 35912 12102 35940 12718
rect 35900 12096 35952 12102
rect 35900 12038 35952 12044
rect 35716 11688 35768 11694
rect 35716 11630 35768 11636
rect 35072 11212 35124 11218
rect 35072 11154 35124 11160
rect 34980 11144 35032 11150
rect 34980 11086 35032 11092
rect 34888 11008 34940 11014
rect 34888 10950 34940 10956
rect 34900 10606 34928 10950
rect 34888 10600 34940 10606
rect 34888 10542 34940 10548
rect 34992 10266 35020 11086
rect 36096 10810 36124 12718
rect 36188 12646 36216 12718
rect 36176 12640 36228 12646
rect 36176 12582 36228 12588
rect 36188 12306 36216 12582
rect 36176 12300 36228 12306
rect 36176 12242 36228 12248
rect 36268 11212 36320 11218
rect 36268 11154 36320 11160
rect 36084 10804 36136 10810
rect 36084 10746 36136 10752
rect 34980 10260 35032 10266
rect 34980 10202 35032 10208
rect 34152 10124 34204 10130
rect 34152 10066 34204 10072
rect 34992 9568 35020 10202
rect 35624 10056 35676 10062
rect 35624 9998 35676 10004
rect 34992 9540 35112 9568
rect 33968 9444 34020 9450
rect 33968 9386 34020 9392
rect 34980 9444 35032 9450
rect 34980 9386 35032 9392
rect 34796 9376 34848 9382
rect 34796 9318 34848 9324
rect 34808 8838 34836 9318
rect 34888 9036 34940 9042
rect 34888 8978 34940 8984
rect 34796 8832 34848 8838
rect 34796 8774 34848 8780
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 33876 8492 33928 8498
rect 33876 8434 33928 8440
rect 33784 8424 33836 8430
rect 33784 8366 33836 8372
rect 33232 8016 33284 8022
rect 33232 7958 33284 7964
rect 33416 8016 33468 8022
rect 33416 7958 33468 7964
rect 33244 7342 33272 7958
rect 33796 7886 33824 8366
rect 33784 7880 33836 7886
rect 33784 7822 33836 7828
rect 33600 7812 33652 7818
rect 33600 7754 33652 7760
rect 33612 7410 33640 7754
rect 33796 7410 33824 7822
rect 33600 7404 33652 7410
rect 33600 7346 33652 7352
rect 33784 7404 33836 7410
rect 33784 7346 33836 7352
rect 33232 7336 33284 7342
rect 33232 7278 33284 7284
rect 33784 7200 33836 7206
rect 33784 7142 33836 7148
rect 33796 6866 33824 7142
rect 33416 6860 33468 6866
rect 33416 6802 33468 6808
rect 33784 6860 33836 6866
rect 33784 6802 33836 6808
rect 33324 6724 33376 6730
rect 33324 6666 33376 6672
rect 33232 6656 33284 6662
rect 33232 6598 33284 6604
rect 33244 6458 33272 6598
rect 33232 6452 33284 6458
rect 33232 6394 33284 6400
rect 33336 6322 33364 6666
rect 33324 6316 33376 6322
rect 33324 6258 33376 6264
rect 33232 5704 33284 5710
rect 33232 5646 33284 5652
rect 33140 4820 33192 4826
rect 33140 4762 33192 4768
rect 33048 4276 33100 4282
rect 33048 4218 33100 4224
rect 32954 4176 33010 4185
rect 32954 4111 33010 4120
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 32956 3392 33008 3398
rect 32956 3334 33008 3340
rect 32968 2990 32996 3334
rect 32956 2984 33008 2990
rect 32956 2926 33008 2932
rect 33060 2854 33088 3470
rect 33244 3194 33272 5646
rect 33324 5160 33376 5166
rect 33324 5102 33376 5108
rect 33336 4486 33364 5102
rect 33428 5030 33456 6802
rect 34072 6254 34100 8570
rect 34520 8492 34572 8498
rect 34520 8434 34572 8440
rect 34532 7954 34560 8434
rect 34900 8430 34928 8978
rect 34888 8424 34940 8430
rect 34888 8366 34940 8372
rect 34900 7954 34928 8366
rect 34992 7954 35020 9386
rect 35084 8974 35112 9540
rect 35348 9512 35400 9518
rect 35348 9454 35400 9460
rect 35440 9512 35492 9518
rect 35440 9454 35492 9460
rect 35072 8968 35124 8974
rect 35072 8910 35124 8916
rect 34520 7948 34572 7954
rect 34520 7890 34572 7896
rect 34888 7948 34940 7954
rect 34888 7890 34940 7896
rect 34980 7948 35032 7954
rect 34980 7890 35032 7896
rect 34336 7336 34388 7342
rect 34336 7278 34388 7284
rect 34060 6248 34112 6254
rect 34060 6190 34112 6196
rect 34244 6248 34296 6254
rect 34244 6190 34296 6196
rect 34072 5710 34100 6190
rect 34060 5704 34112 5710
rect 34060 5646 34112 5652
rect 34256 5030 34284 6190
rect 34348 5710 34376 7278
rect 34900 6866 34928 7890
rect 35360 7274 35388 9454
rect 35452 8430 35480 9454
rect 35636 9110 35664 9998
rect 36280 9654 36308 11154
rect 36372 10266 36400 13194
rect 36544 12776 36596 12782
rect 36544 12718 36596 12724
rect 36452 12232 36504 12238
rect 36452 12174 36504 12180
rect 36464 11694 36492 12174
rect 36452 11688 36504 11694
rect 36452 11630 36504 11636
rect 36464 11014 36492 11630
rect 36556 11218 36584 12718
rect 36648 12374 36676 14894
rect 37188 14544 37240 14550
rect 37188 14486 37240 14492
rect 36820 13864 36872 13870
rect 36820 13806 36872 13812
rect 36832 13462 36860 13806
rect 36820 13456 36872 13462
rect 36820 13398 36872 13404
rect 36636 12368 36688 12374
rect 36636 12310 36688 12316
rect 37200 12102 37228 14486
rect 37384 14006 37412 14962
rect 37648 14408 37700 14414
rect 37648 14350 37700 14356
rect 37660 14006 37688 14350
rect 37372 14000 37424 14006
rect 37372 13942 37424 13948
rect 37648 14000 37700 14006
rect 37648 13942 37700 13948
rect 37384 13734 37412 13942
rect 37372 13728 37424 13734
rect 37372 13670 37424 13676
rect 37752 13462 37780 15506
rect 37740 13456 37792 13462
rect 37740 13398 37792 13404
rect 37464 12776 37516 12782
rect 37464 12718 37516 12724
rect 37370 12472 37426 12481
rect 37370 12407 37426 12416
rect 36728 12096 36780 12102
rect 36728 12038 36780 12044
rect 37188 12096 37240 12102
rect 37188 12038 37240 12044
rect 36740 11694 36768 12038
rect 37384 11830 37412 12407
rect 37372 11824 37424 11830
rect 37372 11766 37424 11772
rect 36636 11688 36688 11694
rect 36636 11630 36688 11636
rect 36728 11688 36780 11694
rect 36728 11630 36780 11636
rect 37096 11688 37148 11694
rect 37148 11648 37228 11676
rect 37096 11630 37148 11636
rect 36544 11212 36596 11218
rect 36544 11154 36596 11160
rect 36648 11082 36676 11630
rect 36820 11212 36872 11218
rect 36820 11154 36872 11160
rect 36636 11076 36688 11082
rect 36636 11018 36688 11024
rect 36452 11008 36504 11014
rect 36452 10950 36504 10956
rect 36360 10260 36412 10266
rect 36360 10202 36412 10208
rect 36268 9648 36320 9654
rect 36268 9590 36320 9596
rect 35900 9512 35952 9518
rect 35900 9454 35952 9460
rect 36452 9512 36504 9518
rect 36452 9454 36504 9460
rect 36728 9512 36780 9518
rect 36728 9454 36780 9460
rect 35624 9104 35676 9110
rect 35624 9046 35676 9052
rect 35440 8424 35492 8430
rect 35440 8366 35492 8372
rect 35716 8424 35768 8430
rect 35716 8366 35768 8372
rect 35348 7268 35400 7274
rect 35348 7210 35400 7216
rect 35452 7206 35480 8366
rect 35624 8356 35676 8362
rect 35544 8316 35624 8344
rect 35544 7342 35572 8316
rect 35624 8298 35676 8304
rect 35532 7336 35584 7342
rect 35532 7278 35584 7284
rect 35440 7200 35492 7206
rect 35440 7142 35492 7148
rect 35544 6866 35572 7278
rect 35728 7041 35756 8366
rect 35912 7936 35940 9454
rect 36084 9036 36136 9042
rect 36084 8978 36136 8984
rect 36096 8634 36124 8978
rect 36084 8628 36136 8634
rect 36084 8570 36136 8576
rect 36176 8356 36228 8362
rect 36176 8298 36228 8304
rect 36084 7948 36136 7954
rect 35912 7908 36084 7936
rect 35714 7032 35770 7041
rect 35714 6967 35770 6976
rect 34888 6860 34940 6866
rect 34888 6802 34940 6808
rect 35532 6860 35584 6866
rect 35532 6802 35584 6808
rect 35912 6186 35940 7908
rect 36188 7936 36216 8298
rect 36464 8242 36492 9454
rect 36636 9444 36688 9450
rect 36636 9386 36688 9392
rect 36648 9178 36676 9386
rect 36740 9178 36768 9454
rect 36832 9382 36860 11154
rect 36912 9920 36964 9926
rect 36912 9862 36964 9868
rect 36820 9376 36872 9382
rect 36820 9318 36872 9324
rect 36636 9172 36688 9178
rect 36636 9114 36688 9120
rect 36728 9172 36780 9178
rect 36728 9114 36780 9120
rect 36832 9042 36860 9318
rect 36820 9036 36872 9042
rect 36820 8978 36872 8984
rect 36728 8968 36780 8974
rect 36728 8910 36780 8916
rect 36544 8560 36596 8566
rect 36544 8502 36596 8508
rect 36556 8412 36584 8502
rect 36740 8412 36768 8910
rect 36556 8384 36768 8412
rect 36820 8424 36872 8430
rect 36820 8366 36872 8372
rect 36464 8214 36676 8242
rect 36268 7948 36320 7954
rect 36188 7908 36268 7936
rect 36084 7890 36136 7896
rect 36268 7890 36320 7896
rect 36360 7404 36412 7410
rect 36360 7346 36412 7352
rect 36084 7336 36136 7342
rect 36084 7278 36136 7284
rect 36176 7336 36228 7342
rect 36176 7278 36228 7284
rect 35990 7168 36046 7177
rect 35990 7103 36046 7112
rect 36004 6866 36032 7103
rect 35992 6860 36044 6866
rect 35992 6802 36044 6808
rect 36004 6390 36032 6802
rect 35992 6384 36044 6390
rect 35992 6326 36044 6332
rect 35900 6180 35952 6186
rect 35900 6122 35952 6128
rect 35072 6112 35124 6118
rect 35072 6054 35124 6060
rect 35084 5914 35112 6054
rect 35072 5908 35124 5914
rect 35072 5850 35124 5856
rect 34612 5840 34664 5846
rect 34612 5782 34664 5788
rect 34336 5704 34388 5710
rect 34388 5652 34560 5658
rect 34336 5646 34560 5652
rect 34348 5642 34560 5646
rect 34348 5636 34572 5642
rect 34348 5630 34520 5636
rect 33416 5024 33468 5030
rect 33416 4966 33468 4972
rect 34244 5024 34296 5030
rect 34244 4966 34296 4972
rect 33324 4480 33376 4486
rect 33324 4422 33376 4428
rect 34242 3224 34298 3233
rect 33232 3188 33284 3194
rect 33232 3130 33284 3136
rect 33324 3188 33376 3194
rect 34242 3159 34298 3168
rect 33324 3130 33376 3136
rect 33048 2848 33100 2854
rect 33048 2790 33100 2796
rect 32864 2304 32916 2310
rect 32864 2246 32916 2252
rect 32772 1896 32824 1902
rect 32772 1838 32824 1844
rect 31404 870 31616 898
rect 31588 800 31616 870
rect 32416 870 32536 898
rect 32416 800 32444 870
rect 33336 800 33364 3130
rect 33966 2680 34022 2689
rect 33966 2615 34022 2624
rect 33980 2582 34008 2615
rect 33968 2576 34020 2582
rect 33968 2518 34020 2524
rect 34256 898 34284 3159
rect 34348 3058 34376 5630
rect 34520 5578 34572 5584
rect 34428 3936 34480 3942
rect 34428 3878 34480 3884
rect 34440 3602 34468 3878
rect 34624 3670 34652 5782
rect 34796 5160 34848 5166
rect 34796 5102 34848 5108
rect 34612 3664 34664 3670
rect 34612 3606 34664 3612
rect 34702 3632 34758 3641
rect 34428 3596 34480 3602
rect 34702 3567 34758 3576
rect 34428 3538 34480 3544
rect 34716 3369 34744 3567
rect 34518 3360 34574 3369
rect 34518 3295 34574 3304
rect 34702 3360 34758 3369
rect 34702 3295 34758 3304
rect 34336 3052 34388 3058
rect 34336 2994 34388 3000
rect 34532 2825 34560 3295
rect 34612 3052 34664 3058
rect 34612 2994 34664 3000
rect 34518 2816 34574 2825
rect 34518 2751 34574 2760
rect 34624 2446 34652 2994
rect 34612 2440 34664 2446
rect 34612 2382 34664 2388
rect 34808 1902 34836 5102
rect 34888 5024 34940 5030
rect 34888 4966 34940 4972
rect 34900 3126 34928 4966
rect 36096 4622 36124 7278
rect 36188 6866 36216 7278
rect 36372 6866 36400 7346
rect 36176 6860 36228 6866
rect 36176 6802 36228 6808
rect 36360 6860 36412 6866
rect 36360 6802 36412 6808
rect 36452 6860 36504 6866
rect 36452 6802 36504 6808
rect 36188 6458 36216 6802
rect 36464 6746 36492 6802
rect 36280 6718 36492 6746
rect 36176 6452 36228 6458
rect 36176 6394 36228 6400
rect 36176 5636 36228 5642
rect 36176 5578 36228 5584
rect 36188 5030 36216 5578
rect 36280 5574 36308 6718
rect 36452 6384 36504 6390
rect 36452 6326 36504 6332
rect 36464 6254 36492 6326
rect 36452 6248 36504 6254
rect 36504 6208 36584 6236
rect 36452 6190 36504 6196
rect 36360 6180 36412 6186
rect 36360 6122 36412 6128
rect 36372 5642 36400 6122
rect 36452 6112 36504 6118
rect 36452 6054 36504 6060
rect 36360 5636 36412 5642
rect 36360 5578 36412 5584
rect 36268 5568 36320 5574
rect 36268 5510 36320 5516
rect 36464 5166 36492 6054
rect 36556 5166 36584 6208
rect 36452 5160 36504 5166
rect 36452 5102 36504 5108
rect 36544 5160 36596 5166
rect 36544 5102 36596 5108
rect 36176 5024 36228 5030
rect 36648 4978 36676 8214
rect 36832 6390 36860 8366
rect 36924 6458 36952 9862
rect 37096 9648 37148 9654
rect 37096 9590 37148 9596
rect 37108 9110 37136 9590
rect 37096 9104 37148 9110
rect 37096 9046 37148 9052
rect 37004 8900 37056 8906
rect 37004 8842 37056 8848
rect 37016 8566 37044 8842
rect 37004 8560 37056 8566
rect 37004 8502 37056 8508
rect 37096 7744 37148 7750
rect 37096 7686 37148 7692
rect 37108 7342 37136 7686
rect 37004 7336 37056 7342
rect 37004 7278 37056 7284
rect 37096 7336 37148 7342
rect 37096 7278 37148 7284
rect 37016 6866 37044 7278
rect 37200 7002 37228 11648
rect 37476 11540 37504 12718
rect 37844 12238 37872 16050
rect 38384 16040 38436 16046
rect 38384 15982 38436 15988
rect 38200 15972 38252 15978
rect 38200 15914 38252 15920
rect 38212 13802 38240 15914
rect 38396 15706 38424 15982
rect 38384 15700 38436 15706
rect 38384 15642 38436 15648
rect 38396 15570 38424 15642
rect 38384 15564 38436 15570
rect 38384 15506 38436 15512
rect 38764 15366 38792 17070
rect 38948 16046 38976 17138
rect 39224 16998 39252 18835
rect 41156 17338 41184 18835
rect 40500 17332 40552 17338
rect 40500 17274 40552 17280
rect 41144 17332 41196 17338
rect 41144 17274 41196 17280
rect 39212 16992 39264 16998
rect 39212 16934 39264 16940
rect 39224 16794 39252 16934
rect 39212 16788 39264 16794
rect 39212 16730 39264 16736
rect 40512 16658 40540 17274
rect 41681 16892 41977 16912
rect 41737 16890 41761 16892
rect 41817 16890 41841 16892
rect 41897 16890 41921 16892
rect 41759 16838 41761 16890
rect 41823 16838 41835 16890
rect 41897 16838 41899 16890
rect 41737 16836 41761 16838
rect 41817 16836 41841 16838
rect 41897 16836 41921 16838
rect 41681 16816 41977 16836
rect 39212 16652 39264 16658
rect 39212 16594 39264 16600
rect 40500 16652 40552 16658
rect 40500 16594 40552 16600
rect 42892 16652 42944 16658
rect 42892 16594 42944 16600
rect 39224 16250 39252 16594
rect 40592 16448 40644 16454
rect 40592 16390 40644 16396
rect 39212 16244 39264 16250
rect 39212 16186 39264 16192
rect 38936 16040 38988 16046
rect 38936 15982 38988 15988
rect 40604 15638 40632 16390
rect 42064 16040 42116 16046
rect 42064 15982 42116 15988
rect 41681 15804 41977 15824
rect 41737 15802 41761 15804
rect 41817 15802 41841 15804
rect 41897 15802 41921 15804
rect 41759 15750 41761 15802
rect 41823 15750 41835 15802
rect 41897 15750 41899 15802
rect 41737 15748 41761 15750
rect 41817 15748 41841 15750
rect 41897 15748 41921 15750
rect 41681 15728 41977 15748
rect 40592 15632 40644 15638
rect 40592 15574 40644 15580
rect 39028 15564 39080 15570
rect 39028 15506 39080 15512
rect 38752 15360 38804 15366
rect 38752 15302 38804 15308
rect 38660 14952 38712 14958
rect 38660 14894 38712 14900
rect 38568 14476 38620 14482
rect 38568 14418 38620 14424
rect 38476 14408 38528 14414
rect 38476 14350 38528 14356
rect 38200 13796 38252 13802
rect 38200 13738 38252 13744
rect 38488 13734 38516 14350
rect 38580 14074 38608 14418
rect 38672 14346 38700 14894
rect 39040 14550 39068 15506
rect 42076 15434 42104 15982
rect 42064 15428 42116 15434
rect 42064 15370 42116 15376
rect 41604 14952 41656 14958
rect 41604 14894 41656 14900
rect 40960 14884 41012 14890
rect 40960 14826 41012 14832
rect 39120 14816 39172 14822
rect 39120 14758 39172 14764
rect 39132 14618 39160 14758
rect 39120 14612 39172 14618
rect 39120 14554 39172 14560
rect 39028 14544 39080 14550
rect 39028 14486 39080 14492
rect 39856 14408 39908 14414
rect 39856 14350 39908 14356
rect 38660 14340 38712 14346
rect 38660 14282 38712 14288
rect 39396 14340 39448 14346
rect 39396 14282 39448 14288
rect 38568 14068 38620 14074
rect 38568 14010 38620 14016
rect 38476 13728 38528 13734
rect 38476 13670 38528 13676
rect 38488 13394 38516 13670
rect 38384 13388 38436 13394
rect 38384 13330 38436 13336
rect 38476 13388 38528 13394
rect 38476 13330 38528 13336
rect 38396 12850 38424 13330
rect 38384 12844 38436 12850
rect 38384 12786 38436 12792
rect 37832 12232 37884 12238
rect 37832 12174 37884 12180
rect 37648 11552 37700 11558
rect 37476 11512 37648 11540
rect 37648 11494 37700 11500
rect 37740 10124 37792 10130
rect 37740 10066 37792 10072
rect 37278 9616 37334 9625
rect 37278 9551 37280 9560
rect 37332 9551 37334 9560
rect 37280 9522 37332 9528
rect 37280 9444 37332 9450
rect 37280 9386 37332 9392
rect 37292 8430 37320 9386
rect 37752 8838 37780 10066
rect 37924 8900 37976 8906
rect 37924 8842 37976 8848
rect 37740 8832 37792 8838
rect 37740 8774 37792 8780
rect 37280 8424 37332 8430
rect 37280 8366 37332 8372
rect 37372 8016 37424 8022
rect 37372 7958 37424 7964
rect 37280 7268 37332 7274
rect 37280 7210 37332 7216
rect 37188 6996 37240 7002
rect 37188 6938 37240 6944
rect 37004 6860 37056 6866
rect 37004 6802 37056 6808
rect 36912 6452 36964 6458
rect 36912 6394 36964 6400
rect 36820 6384 36872 6390
rect 36820 6326 36872 6332
rect 36728 5364 36780 5370
rect 36728 5306 36780 5312
rect 36740 5166 36768 5306
rect 36728 5160 36780 5166
rect 36728 5102 36780 5108
rect 36176 4966 36228 4972
rect 36556 4950 36676 4978
rect 36360 4684 36412 4690
rect 36360 4626 36412 4632
rect 36084 4616 36136 4622
rect 35346 4584 35402 4593
rect 36084 4558 36136 4564
rect 35346 4519 35348 4528
rect 35400 4519 35402 4528
rect 35348 4490 35400 4496
rect 34980 4480 35032 4486
rect 34980 4422 35032 4428
rect 34992 4214 35020 4422
rect 34980 4208 35032 4214
rect 34980 4150 35032 4156
rect 34992 4078 35020 4150
rect 34980 4072 35032 4078
rect 34980 4014 35032 4020
rect 36084 4072 36136 4078
rect 36084 4014 36136 4020
rect 35716 3936 35768 3942
rect 35716 3878 35768 3884
rect 34978 3632 35034 3641
rect 34978 3567 35034 3576
rect 34888 3120 34940 3126
rect 34888 3062 34940 3068
rect 34796 1896 34848 1902
rect 34796 1838 34848 1844
rect 34164 870 34284 898
rect 34164 800 34192 870
rect 34992 800 35020 3567
rect 35532 3528 35584 3534
rect 35530 3496 35532 3505
rect 35584 3496 35586 3505
rect 35530 3431 35586 3440
rect 35728 2990 35756 3878
rect 35992 3120 36044 3126
rect 35992 3062 36044 3068
rect 35624 2984 35676 2990
rect 35624 2926 35676 2932
rect 35716 2984 35768 2990
rect 35716 2926 35768 2932
rect 35636 2802 35664 2926
rect 36004 2854 36032 3062
rect 35992 2848 36044 2854
rect 35636 2774 35940 2802
rect 35992 2790 36044 2796
rect 35912 2514 35940 2774
rect 35900 2508 35952 2514
rect 35900 2450 35952 2456
rect 35912 800 35940 2450
rect 36096 2446 36124 4014
rect 36176 3936 36228 3942
rect 36176 3878 36228 3884
rect 36188 3670 36216 3878
rect 36266 3768 36322 3777
rect 36266 3703 36322 3712
rect 36280 3670 36308 3703
rect 36176 3664 36228 3670
rect 36176 3606 36228 3612
rect 36268 3664 36320 3670
rect 36268 3606 36320 3612
rect 36188 2689 36216 3606
rect 36372 3534 36400 4626
rect 36360 3528 36412 3534
rect 36360 3470 36412 3476
rect 36268 2916 36320 2922
rect 36268 2858 36320 2864
rect 36174 2680 36230 2689
rect 36174 2615 36230 2624
rect 36280 2514 36308 2858
rect 36268 2508 36320 2514
rect 36268 2450 36320 2456
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 36096 1834 36124 2382
rect 36280 2038 36308 2450
rect 36268 2032 36320 2038
rect 36268 1974 36320 1980
rect 36372 1970 36400 3470
rect 36556 2825 36584 4950
rect 36636 4004 36688 4010
rect 36636 3946 36688 3952
rect 36648 3126 36676 3946
rect 36832 3913 36860 6326
rect 36924 6254 36952 6394
rect 36912 6248 36964 6254
rect 36912 6190 36964 6196
rect 37096 6248 37148 6254
rect 37096 6190 37148 6196
rect 37108 5166 37136 6190
rect 37200 5930 37228 6938
rect 37292 6769 37320 7210
rect 37278 6760 37334 6769
rect 37278 6695 37334 6704
rect 37200 5902 37320 5930
rect 37188 5772 37240 5778
rect 37188 5714 37240 5720
rect 37200 5166 37228 5714
rect 37292 5574 37320 5902
rect 37280 5568 37332 5574
rect 37280 5510 37332 5516
rect 36912 5160 36964 5166
rect 36912 5102 36964 5108
rect 37096 5160 37148 5166
rect 37096 5102 37148 5108
rect 37188 5160 37240 5166
rect 37188 5102 37240 5108
rect 36924 5030 36952 5102
rect 36912 5024 36964 5030
rect 36912 4966 36964 4972
rect 37200 4758 37228 5102
rect 37188 4752 37240 4758
rect 37188 4694 37240 4700
rect 36818 3904 36874 3913
rect 36818 3839 36874 3848
rect 37200 3602 37228 4694
rect 37280 4616 37332 4622
rect 37280 4558 37332 4564
rect 37292 4078 37320 4558
rect 37384 4282 37412 7958
rect 37752 7954 37780 8774
rect 37740 7948 37792 7954
rect 37740 7890 37792 7896
rect 37752 7002 37780 7890
rect 37740 6996 37792 7002
rect 37740 6938 37792 6944
rect 37556 6860 37608 6866
rect 37556 6802 37608 6808
rect 37740 6860 37792 6866
rect 37740 6802 37792 6808
rect 37568 6236 37596 6802
rect 37648 6248 37700 6254
rect 37568 6208 37648 6236
rect 37648 6190 37700 6196
rect 37464 4480 37516 4486
rect 37464 4422 37516 4428
rect 37372 4276 37424 4282
rect 37372 4218 37424 4224
rect 37476 4146 37504 4422
rect 37464 4140 37516 4146
rect 37464 4082 37516 4088
rect 37280 4072 37332 4078
rect 37280 4014 37332 4020
rect 36728 3596 36780 3602
rect 36728 3538 36780 3544
rect 37188 3596 37240 3602
rect 37188 3538 37240 3544
rect 36636 3120 36688 3126
rect 36636 3062 36688 3068
rect 36740 3058 36768 3538
rect 37660 3398 37688 6190
rect 37752 4214 37780 6802
rect 37936 5914 37964 8842
rect 38292 8424 38344 8430
rect 38292 8366 38344 8372
rect 38016 7744 38068 7750
rect 38016 7686 38068 7692
rect 37924 5908 37976 5914
rect 37924 5850 37976 5856
rect 38028 5370 38056 7686
rect 38108 7404 38160 7410
rect 38108 7346 38160 7352
rect 38016 5364 38068 5370
rect 38016 5306 38068 5312
rect 38120 4758 38148 7346
rect 38200 6860 38252 6866
rect 38304 6848 38332 8366
rect 38580 7410 38608 14010
rect 38672 13870 38700 14282
rect 39120 14272 39172 14278
rect 39120 14214 39172 14220
rect 39132 13938 39160 14214
rect 39120 13932 39172 13938
rect 39120 13874 39172 13880
rect 39408 13870 39436 14282
rect 39868 13870 39896 14350
rect 40776 14340 40828 14346
rect 40776 14282 40828 14288
rect 38660 13864 38712 13870
rect 38660 13806 38712 13812
rect 38844 13864 38896 13870
rect 38844 13806 38896 13812
rect 39396 13864 39448 13870
rect 39396 13806 39448 13812
rect 39856 13864 39908 13870
rect 39856 13806 39908 13812
rect 38856 12782 38884 13806
rect 39408 13394 39436 13806
rect 39396 13388 39448 13394
rect 39396 13330 39448 13336
rect 40500 13184 40552 13190
rect 40500 13126 40552 13132
rect 40512 12850 40540 13126
rect 40788 12986 40816 14282
rect 40592 12980 40644 12986
rect 40592 12922 40644 12928
rect 40776 12980 40828 12986
rect 40776 12922 40828 12928
rect 40604 12866 40632 12922
rect 40500 12844 40552 12850
rect 40604 12838 40816 12866
rect 40500 12786 40552 12792
rect 38844 12776 38896 12782
rect 38844 12718 38896 12724
rect 38752 12232 38804 12238
rect 38752 12174 38804 12180
rect 39028 12232 39080 12238
rect 39028 12174 39080 12180
rect 38764 11150 38792 12174
rect 38936 11892 38988 11898
rect 38936 11834 38988 11840
rect 38752 11144 38804 11150
rect 38752 11086 38804 11092
rect 38844 11076 38896 11082
rect 38844 11018 38896 11024
rect 38856 10606 38884 11018
rect 38948 10606 38976 11834
rect 39040 10742 39068 12174
rect 39672 12096 39724 12102
rect 39672 12038 39724 12044
rect 40132 12096 40184 12102
rect 40132 12038 40184 12044
rect 39684 11937 39712 12038
rect 39670 11928 39726 11937
rect 40144 11898 40172 12038
rect 39670 11863 39726 11872
rect 40132 11892 40184 11898
rect 40132 11834 40184 11840
rect 40512 11354 40540 12786
rect 40684 12776 40736 12782
rect 40684 12718 40736 12724
rect 40696 12102 40724 12718
rect 40684 12096 40736 12102
rect 40684 12038 40736 12044
rect 40500 11348 40552 11354
rect 40500 11290 40552 11296
rect 39212 11144 39264 11150
rect 39212 11086 39264 11092
rect 39488 11144 39540 11150
rect 39488 11086 39540 11092
rect 39028 10736 39080 10742
rect 39028 10678 39080 10684
rect 39224 10674 39252 11086
rect 39212 10668 39264 10674
rect 39212 10610 39264 10616
rect 38660 10600 38712 10606
rect 38660 10542 38712 10548
rect 38844 10600 38896 10606
rect 38844 10542 38896 10548
rect 38936 10600 38988 10606
rect 38936 10542 38988 10548
rect 38672 9110 38700 10542
rect 38856 10062 38884 10542
rect 39500 10198 39528 11086
rect 39488 10192 39540 10198
rect 39488 10134 39540 10140
rect 40512 10130 40540 11290
rect 39580 10124 39632 10130
rect 39580 10066 39632 10072
rect 40500 10124 40552 10130
rect 40500 10066 40552 10072
rect 38844 10056 38896 10062
rect 38844 9998 38896 10004
rect 38752 9512 38804 9518
rect 38752 9454 38804 9460
rect 38660 9104 38712 9110
rect 38660 9046 38712 9052
rect 38764 8956 38792 9454
rect 39304 9444 39356 9450
rect 39304 9386 39356 9392
rect 39316 9042 39344 9386
rect 39304 9036 39356 9042
rect 39304 8978 39356 8984
rect 38672 8928 38792 8956
rect 38568 7404 38620 7410
rect 38568 7346 38620 7352
rect 38568 7200 38620 7206
rect 38566 7168 38568 7177
rect 38620 7168 38622 7177
rect 38566 7103 38622 7112
rect 38252 6820 38332 6848
rect 38200 6802 38252 6808
rect 38672 5658 38700 8928
rect 39316 8634 39344 8978
rect 39304 8628 39356 8634
rect 39304 8570 39356 8576
rect 39488 8628 39540 8634
rect 39488 8570 39540 8576
rect 39316 7954 39344 8570
rect 39304 7948 39356 7954
rect 39304 7890 39356 7896
rect 38844 7880 38896 7886
rect 38844 7822 38896 7828
rect 38752 7268 38804 7274
rect 38752 7210 38804 7216
rect 38764 7177 38792 7210
rect 38750 7168 38806 7177
rect 38750 7103 38806 7112
rect 38752 6860 38804 6866
rect 38752 6802 38804 6808
rect 38764 5778 38792 6802
rect 38856 6458 38884 7822
rect 38936 6860 38988 6866
rect 38936 6802 38988 6808
rect 38844 6452 38896 6458
rect 38844 6394 38896 6400
rect 38752 5772 38804 5778
rect 38752 5714 38804 5720
rect 38672 5630 38792 5658
rect 38108 4752 38160 4758
rect 38108 4694 38160 4700
rect 38384 4684 38436 4690
rect 38384 4626 38436 4632
rect 38396 4570 38424 4626
rect 37832 4548 37884 4554
rect 38396 4542 38516 4570
rect 37832 4490 37884 4496
rect 37740 4208 37792 4214
rect 37740 4150 37792 4156
rect 37844 3602 37872 4490
rect 38108 4480 38160 4486
rect 38108 4422 38160 4428
rect 37924 4140 37976 4146
rect 37924 4082 37976 4088
rect 37832 3596 37884 3602
rect 37832 3538 37884 3544
rect 37648 3392 37700 3398
rect 37648 3334 37700 3340
rect 36728 3052 36780 3058
rect 36728 2994 36780 3000
rect 37936 2990 37964 4082
rect 38120 3194 38148 4422
rect 38200 4004 38252 4010
rect 38200 3946 38252 3952
rect 38108 3188 38160 3194
rect 38108 3130 38160 3136
rect 37924 2984 37976 2990
rect 37924 2926 37976 2932
rect 36542 2816 36598 2825
rect 36542 2751 36598 2760
rect 37936 2514 37964 2926
rect 38120 2582 38148 3130
rect 38212 3058 38240 3946
rect 38488 3534 38516 4542
rect 38660 4480 38712 4486
rect 38660 4422 38712 4428
rect 38568 4140 38620 4146
rect 38568 4082 38620 4088
rect 38476 3528 38528 3534
rect 38476 3470 38528 3476
rect 38200 3052 38252 3058
rect 38200 2994 38252 3000
rect 38488 2990 38516 3470
rect 38580 3466 38608 4082
rect 38568 3460 38620 3466
rect 38568 3402 38620 3408
rect 38476 2984 38528 2990
rect 38476 2926 38528 2932
rect 38108 2576 38160 2582
rect 38108 2518 38160 2524
rect 38672 2514 38700 4422
rect 38764 2961 38792 5630
rect 38856 3670 38884 6394
rect 38948 6390 38976 6802
rect 38936 6384 38988 6390
rect 38936 6326 38988 6332
rect 39120 6248 39172 6254
rect 39120 6190 39172 6196
rect 39028 5908 39080 5914
rect 39028 5850 39080 5856
rect 39040 5166 39068 5850
rect 39132 5846 39160 6190
rect 39120 5840 39172 5846
rect 39120 5782 39172 5788
rect 39028 5160 39080 5166
rect 39028 5102 39080 5108
rect 39120 5160 39172 5166
rect 39120 5102 39172 5108
rect 38936 5092 38988 5098
rect 38936 5034 38988 5040
rect 38948 4690 38976 5034
rect 38936 4684 38988 4690
rect 38936 4626 38988 4632
rect 38948 4146 38976 4626
rect 38936 4140 38988 4146
rect 38936 4082 38988 4088
rect 38844 3664 38896 3670
rect 38844 3606 38896 3612
rect 39028 3596 39080 3602
rect 39028 3538 39080 3544
rect 39040 3505 39068 3538
rect 39026 3496 39082 3505
rect 39026 3431 39082 3440
rect 39132 3058 39160 5102
rect 39316 4078 39344 7890
rect 39500 6662 39528 8570
rect 39592 8022 39620 10066
rect 39948 9376 40000 9382
rect 39948 9318 40000 9324
rect 39960 9042 39988 9318
rect 39948 9036 40000 9042
rect 39948 8978 40000 8984
rect 40040 8832 40092 8838
rect 40040 8774 40092 8780
rect 40052 8430 40080 8774
rect 40040 8424 40092 8430
rect 40040 8366 40092 8372
rect 39764 8288 39816 8294
rect 39764 8230 39816 8236
rect 40684 8288 40736 8294
rect 40684 8230 40736 8236
rect 39776 8090 39804 8230
rect 39764 8084 39816 8090
rect 39764 8026 39816 8032
rect 39580 8016 39632 8022
rect 39580 7958 39632 7964
rect 40316 7948 40368 7954
rect 40316 7890 40368 7896
rect 40328 7478 40356 7890
rect 40408 7744 40460 7750
rect 40408 7686 40460 7692
rect 40316 7472 40368 7478
rect 40316 7414 40368 7420
rect 39488 6656 39540 6662
rect 39488 6598 39540 6604
rect 39396 6316 39448 6322
rect 39396 6258 39448 6264
rect 39408 5778 39436 6258
rect 39500 6186 39528 6598
rect 39672 6384 39724 6390
rect 39672 6326 39724 6332
rect 39488 6180 39540 6186
rect 39488 6122 39540 6128
rect 39488 5840 39540 5846
rect 39488 5782 39540 5788
rect 39396 5772 39448 5778
rect 39396 5714 39448 5720
rect 39500 5166 39528 5782
rect 39684 5166 39712 6326
rect 40328 5166 40356 7414
rect 40420 6866 40448 7686
rect 40696 7410 40724 8230
rect 40684 7404 40736 7410
rect 40684 7346 40736 7352
rect 40408 6860 40460 6866
rect 40408 6802 40460 6808
rect 40684 6452 40736 6458
rect 40684 6394 40736 6400
rect 40696 6254 40724 6394
rect 40684 6248 40736 6254
rect 40684 6190 40736 6196
rect 40408 6180 40460 6186
rect 40408 6122 40460 6128
rect 39488 5160 39540 5166
rect 39488 5102 39540 5108
rect 39672 5160 39724 5166
rect 39672 5102 39724 5108
rect 40316 5160 40368 5166
rect 40316 5102 40368 5108
rect 40040 4752 40092 4758
rect 40040 4694 40092 4700
rect 40052 4146 40080 4694
rect 40420 4554 40448 6122
rect 40592 5568 40644 5574
rect 40592 5510 40644 5516
rect 40604 5234 40632 5510
rect 40592 5228 40644 5234
rect 40592 5170 40644 5176
rect 40408 4548 40460 4554
rect 40408 4490 40460 4496
rect 40040 4140 40092 4146
rect 40040 4082 40092 4088
rect 39304 4072 39356 4078
rect 39304 4014 39356 4020
rect 39580 4072 39632 4078
rect 39580 4014 39632 4020
rect 39212 4004 39264 4010
rect 39212 3946 39264 3952
rect 39224 3602 39252 3946
rect 39592 3738 39620 4014
rect 39580 3732 39632 3738
rect 39580 3674 39632 3680
rect 40420 3602 40448 4490
rect 40500 4140 40552 4146
rect 40500 4082 40552 4088
rect 39212 3596 39264 3602
rect 39212 3538 39264 3544
rect 40408 3596 40460 3602
rect 40408 3538 40460 3544
rect 40512 3534 40540 4082
rect 40500 3528 40552 3534
rect 40500 3470 40552 3476
rect 40788 3126 40816 12838
rect 40972 8401 41000 14826
rect 41616 14618 41644 14894
rect 41681 14716 41977 14736
rect 41737 14714 41761 14716
rect 41817 14714 41841 14716
rect 41897 14714 41921 14716
rect 41759 14662 41761 14714
rect 41823 14662 41835 14714
rect 41897 14662 41899 14714
rect 41737 14660 41761 14662
rect 41817 14660 41841 14662
rect 41897 14660 41921 14662
rect 41681 14640 41977 14660
rect 42076 14618 42104 15370
rect 41604 14612 41656 14618
rect 41604 14554 41656 14560
rect 42064 14612 42116 14618
rect 42064 14554 42116 14560
rect 41681 13628 41977 13648
rect 41737 13626 41761 13628
rect 41817 13626 41841 13628
rect 41897 13626 41921 13628
rect 41759 13574 41761 13626
rect 41823 13574 41835 13626
rect 41897 13574 41899 13626
rect 41737 13572 41761 13574
rect 41817 13572 41841 13574
rect 41897 13572 41921 13574
rect 41681 13552 41977 13572
rect 42904 13530 42932 16594
rect 43088 16454 43116 18835
rect 45020 17338 45048 18835
rect 45008 17332 45060 17338
rect 45008 17274 45060 17280
rect 43996 17128 44048 17134
rect 43996 17070 44048 17076
rect 44272 17128 44324 17134
rect 44272 17070 44324 17076
rect 44008 16658 44036 17070
rect 43996 16652 44048 16658
rect 43996 16594 44048 16600
rect 43720 16584 43772 16590
rect 43720 16526 43772 16532
rect 43076 16448 43128 16454
rect 43076 16390 43128 16396
rect 43088 16046 43116 16390
rect 43076 16040 43128 16046
rect 43076 15982 43128 15988
rect 43628 15972 43680 15978
rect 43628 15914 43680 15920
rect 43640 15638 43668 15914
rect 43628 15632 43680 15638
rect 43628 15574 43680 15580
rect 43536 15428 43588 15434
rect 43536 15370 43588 15376
rect 43548 15162 43576 15370
rect 43732 15366 43760 16526
rect 44284 16250 44312 17070
rect 44272 16244 44324 16250
rect 44272 16186 44324 16192
rect 44088 16040 44140 16046
rect 44088 15982 44140 15988
rect 44548 16040 44600 16046
rect 44548 15982 44600 15988
rect 44732 16040 44784 16046
rect 44732 15982 44784 15988
rect 44100 15366 44128 15982
rect 44456 15972 44508 15978
rect 44456 15914 44508 15920
rect 44180 15564 44232 15570
rect 44180 15506 44232 15512
rect 43720 15360 43772 15366
rect 43720 15302 43772 15308
rect 44088 15360 44140 15366
rect 44088 15302 44140 15308
rect 43536 15156 43588 15162
rect 43536 15098 43588 15104
rect 43536 14816 43588 14822
rect 43536 14758 43588 14764
rect 42892 13524 42944 13530
rect 42892 13466 42944 13472
rect 41328 13456 41380 13462
rect 41328 13398 41380 13404
rect 42064 13456 42116 13462
rect 42064 13398 42116 13404
rect 41144 12368 41196 12374
rect 41144 12310 41196 12316
rect 41156 11694 41184 12310
rect 41236 11756 41288 11762
rect 41236 11698 41288 11704
rect 41144 11688 41196 11694
rect 41248 11665 41276 11698
rect 41144 11630 41196 11636
rect 41234 11656 41290 11665
rect 41234 11591 41290 11600
rect 41340 11150 41368 13398
rect 41604 13388 41656 13394
rect 41604 13330 41656 13336
rect 41420 13184 41472 13190
rect 41420 13126 41472 13132
rect 41432 12442 41460 13126
rect 41420 12436 41472 12442
rect 41420 12378 41472 12384
rect 41420 12300 41472 12306
rect 41420 12242 41472 12248
rect 41512 12300 41564 12306
rect 41512 12242 41564 12248
rect 41432 11762 41460 12242
rect 41420 11756 41472 11762
rect 41420 11698 41472 11704
rect 41420 11620 41472 11626
rect 41420 11562 41472 11568
rect 41432 11354 41460 11562
rect 41420 11348 41472 11354
rect 41420 11290 41472 11296
rect 41420 11212 41472 11218
rect 41420 11154 41472 11160
rect 41328 11144 41380 11150
rect 41328 11086 41380 11092
rect 41432 10198 41460 11154
rect 41420 10192 41472 10198
rect 41420 10134 41472 10140
rect 41418 9616 41474 9625
rect 41524 9586 41552 12242
rect 41616 11830 41644 13330
rect 41681 12540 41977 12560
rect 41737 12538 41761 12540
rect 41817 12538 41841 12540
rect 41897 12538 41921 12540
rect 41759 12486 41761 12538
rect 41823 12486 41835 12538
rect 41897 12486 41899 12538
rect 41737 12484 41761 12486
rect 41817 12484 41841 12486
rect 41897 12484 41921 12486
rect 41681 12464 41977 12484
rect 42076 12306 42104 13398
rect 42064 12300 42116 12306
rect 42064 12242 42116 12248
rect 42248 12300 42300 12306
rect 42248 12242 42300 12248
rect 41972 12232 42024 12238
rect 41972 12174 42024 12180
rect 42156 12232 42208 12238
rect 42156 12174 42208 12180
rect 41604 11824 41656 11830
rect 41604 11766 41656 11772
rect 41984 11762 42012 12174
rect 41972 11756 42024 11762
rect 41972 11698 42024 11704
rect 41681 11452 41977 11472
rect 41737 11450 41761 11452
rect 41817 11450 41841 11452
rect 41897 11450 41921 11452
rect 41759 11398 41761 11450
rect 41823 11398 41835 11450
rect 41897 11398 41899 11450
rect 41737 11396 41761 11398
rect 41817 11396 41841 11398
rect 41897 11396 41921 11398
rect 41681 11376 41977 11396
rect 41681 10364 41977 10384
rect 41737 10362 41761 10364
rect 41817 10362 41841 10364
rect 41897 10362 41921 10364
rect 41759 10310 41761 10362
rect 41823 10310 41835 10362
rect 41897 10310 41899 10362
rect 41737 10308 41761 10310
rect 41817 10308 41841 10310
rect 41897 10308 41921 10310
rect 41681 10288 41977 10308
rect 42168 10130 42196 12174
rect 42260 11558 42288 12242
rect 42340 11688 42392 11694
rect 42340 11630 42392 11636
rect 42616 11688 42668 11694
rect 42616 11630 42668 11636
rect 42248 11552 42300 11558
rect 42248 11494 42300 11500
rect 42352 10674 42380 11630
rect 42628 11218 42656 11630
rect 42904 11626 42932 13466
rect 43076 13388 43128 13394
rect 43076 13330 43128 13336
rect 43168 13388 43220 13394
rect 43168 13330 43220 13336
rect 43088 12986 43116 13330
rect 43076 12980 43128 12986
rect 43076 12922 43128 12928
rect 43180 12850 43208 13330
rect 43168 12844 43220 12850
rect 43168 12786 43220 12792
rect 43444 12708 43496 12714
rect 43444 12650 43496 12656
rect 43456 12170 43484 12650
rect 43444 12164 43496 12170
rect 43444 12106 43496 12112
rect 42892 11620 42944 11626
rect 42892 11562 42944 11568
rect 43168 11552 43220 11558
rect 43168 11494 43220 11500
rect 43180 11218 43208 11494
rect 42616 11212 42668 11218
rect 42616 11154 42668 11160
rect 43168 11212 43220 11218
rect 43168 11154 43220 11160
rect 43548 11014 43576 14758
rect 43720 14544 43772 14550
rect 43720 14486 43772 14492
rect 43628 14476 43680 14482
rect 43628 14418 43680 14424
rect 43536 11008 43588 11014
rect 43536 10950 43588 10956
rect 42340 10668 42392 10674
rect 42340 10610 42392 10616
rect 42432 10600 42484 10606
rect 42432 10542 42484 10548
rect 41604 10124 41656 10130
rect 41604 10066 41656 10072
rect 42156 10124 42208 10130
rect 42156 10066 42208 10072
rect 41418 9551 41474 9560
rect 41512 9580 41564 9586
rect 41432 9518 41460 9551
rect 41512 9522 41564 9528
rect 41420 9512 41472 9518
rect 41420 9454 41472 9460
rect 41616 9110 41644 10066
rect 42444 9994 42472 10542
rect 42432 9988 42484 9994
rect 42432 9930 42484 9936
rect 42800 9648 42852 9654
rect 41892 9574 42288 9602
rect 42800 9590 42852 9596
rect 41892 9518 41920 9574
rect 41880 9512 41932 9518
rect 41880 9454 41932 9460
rect 42064 9512 42116 9518
rect 42064 9454 42116 9460
rect 41681 9276 41977 9296
rect 41737 9274 41761 9276
rect 41817 9274 41841 9276
rect 41897 9274 41921 9276
rect 41759 9222 41761 9274
rect 41823 9222 41835 9274
rect 41897 9222 41899 9274
rect 41737 9220 41761 9222
rect 41817 9220 41841 9222
rect 41897 9220 41921 9222
rect 41681 9200 41977 9220
rect 41604 9104 41656 9110
rect 41604 9046 41656 9052
rect 41328 8900 41380 8906
rect 41328 8842 41380 8848
rect 40958 8392 41014 8401
rect 40958 8327 41014 8336
rect 41234 8392 41290 8401
rect 41234 8327 41290 8336
rect 41248 7954 41276 8327
rect 41236 7948 41288 7954
rect 41236 7890 41288 7896
rect 40866 7440 40922 7449
rect 40866 7375 40922 7384
rect 40880 6866 40908 7375
rect 41340 7274 41368 8842
rect 42076 8634 42104 9454
rect 42154 8664 42210 8673
rect 42064 8628 42116 8634
rect 42154 8599 42210 8608
rect 42064 8570 42116 8576
rect 42168 8566 42196 8599
rect 42156 8560 42208 8566
rect 42156 8502 42208 8508
rect 41420 8424 41472 8430
rect 41420 8366 41472 8372
rect 42156 8424 42208 8430
rect 42156 8366 42208 8372
rect 41432 7426 41460 8366
rect 42168 8265 42196 8366
rect 42154 8256 42210 8265
rect 41681 8188 41977 8208
rect 42154 8191 42210 8200
rect 41737 8186 41761 8188
rect 41817 8186 41841 8188
rect 41897 8186 41921 8188
rect 41759 8134 41761 8186
rect 41823 8134 41835 8186
rect 41897 8134 41899 8186
rect 41737 8132 41761 8134
rect 41817 8132 41841 8134
rect 41897 8132 41921 8134
rect 41681 8112 41977 8132
rect 42260 7954 42288 9574
rect 42812 8566 42840 9590
rect 43260 9580 43312 9586
rect 43260 9522 43312 9528
rect 43272 9110 43300 9522
rect 43352 9376 43404 9382
rect 43352 9318 43404 9324
rect 43260 9104 43312 9110
rect 43260 9046 43312 9052
rect 42340 8560 42392 8566
rect 42340 8502 42392 8508
rect 42800 8560 42852 8566
rect 42800 8502 42852 8508
rect 42352 8022 42380 8502
rect 42432 8424 42484 8430
rect 42892 8424 42944 8430
rect 42484 8384 42564 8412
rect 42432 8366 42484 8372
rect 42340 8016 42392 8022
rect 42340 7958 42392 7964
rect 41604 7948 41656 7954
rect 41604 7890 41656 7896
rect 42248 7948 42300 7954
rect 42248 7890 42300 7896
rect 41432 7398 41552 7426
rect 41328 7268 41380 7274
rect 41328 7210 41380 7216
rect 41234 7032 41290 7041
rect 41234 6967 41290 6976
rect 41248 6934 41276 6967
rect 41236 6928 41288 6934
rect 41236 6870 41288 6876
rect 40868 6860 40920 6866
rect 40868 6802 40920 6808
rect 41052 6724 41104 6730
rect 41052 6666 41104 6672
rect 40868 5772 40920 5778
rect 40868 5714 40920 5720
rect 40880 5370 40908 5714
rect 40868 5364 40920 5370
rect 40868 5306 40920 5312
rect 40960 5364 41012 5370
rect 40960 5306 41012 5312
rect 40972 5234 41000 5306
rect 40960 5228 41012 5234
rect 40960 5170 41012 5176
rect 40868 4616 40920 4622
rect 40868 4558 40920 4564
rect 40880 4146 40908 4558
rect 41064 4282 41092 6666
rect 41236 4616 41288 4622
rect 41236 4558 41288 4564
rect 41052 4276 41104 4282
rect 41052 4218 41104 4224
rect 40868 4140 40920 4146
rect 40868 4082 40920 4088
rect 41248 3942 41276 4558
rect 41144 3936 41196 3942
rect 41144 3878 41196 3884
rect 41236 3936 41288 3942
rect 41236 3878 41288 3884
rect 41156 3466 41184 3878
rect 41144 3460 41196 3466
rect 41144 3402 41196 3408
rect 41248 3398 41276 3878
rect 41236 3392 41288 3398
rect 41340 3369 41368 7210
rect 41524 6882 41552 7398
rect 41432 6854 41552 6882
rect 41432 6254 41460 6854
rect 41616 6798 41644 7890
rect 42156 7812 42208 7818
rect 42352 7800 42380 7958
rect 42208 7772 42380 7800
rect 42156 7754 42208 7760
rect 42156 7336 42208 7342
rect 42156 7278 42208 7284
rect 42168 7206 42196 7278
rect 42156 7200 42208 7206
rect 42156 7142 42208 7148
rect 41681 7100 41977 7120
rect 41737 7098 41761 7100
rect 41817 7098 41841 7100
rect 41897 7098 41921 7100
rect 41759 7046 41761 7098
rect 41823 7046 41835 7098
rect 41897 7046 41899 7098
rect 41737 7044 41761 7046
rect 41817 7044 41841 7046
rect 41897 7044 41921 7046
rect 41681 7024 41977 7044
rect 41972 6860 42024 6866
rect 41972 6802 42024 6808
rect 41604 6792 41656 6798
rect 41604 6734 41656 6740
rect 41694 6488 41750 6497
rect 41984 6458 42012 6802
rect 41694 6423 41750 6432
rect 41972 6452 42024 6458
rect 41708 6322 41736 6423
rect 41972 6394 42024 6400
rect 42168 6361 42196 7142
rect 42536 6848 42564 8384
rect 42892 8366 42944 8372
rect 42904 7410 42932 8366
rect 42892 7404 42944 7410
rect 42892 7346 42944 7352
rect 43076 7336 43128 7342
rect 43076 7278 43128 7284
rect 42708 6860 42760 6866
rect 42536 6820 42708 6848
rect 42708 6802 42760 6808
rect 42616 6656 42668 6662
rect 42616 6598 42668 6604
rect 42340 6452 42392 6458
rect 42340 6394 42392 6400
rect 42154 6352 42210 6361
rect 41696 6316 41748 6322
rect 42154 6287 42210 6296
rect 41696 6258 41748 6264
rect 41420 6248 41472 6254
rect 41420 6190 41472 6196
rect 42248 6248 42300 6254
rect 42248 6190 42300 6196
rect 41681 6012 41977 6032
rect 41737 6010 41761 6012
rect 41817 6010 41841 6012
rect 41897 6010 41921 6012
rect 41759 5958 41761 6010
rect 41823 5958 41835 6010
rect 41897 5958 41899 6010
rect 41737 5956 41761 5958
rect 41817 5956 41841 5958
rect 41897 5956 41921 5958
rect 41681 5936 41977 5956
rect 42064 5568 42116 5574
rect 42064 5510 42116 5516
rect 41418 5264 41474 5273
rect 41418 5199 41474 5208
rect 41604 5228 41656 5234
rect 41432 5166 41460 5199
rect 41604 5170 41656 5176
rect 41420 5160 41472 5166
rect 41420 5102 41472 5108
rect 41616 3738 41644 5170
rect 41681 4924 41977 4944
rect 41737 4922 41761 4924
rect 41817 4922 41841 4924
rect 41897 4922 41921 4924
rect 41759 4870 41761 4922
rect 41823 4870 41835 4922
rect 41897 4870 41899 4922
rect 41737 4868 41761 4870
rect 41817 4868 41841 4870
rect 41897 4868 41921 4870
rect 41681 4848 41977 4868
rect 42076 4706 42104 5510
rect 42260 5166 42288 6190
rect 42352 6186 42380 6394
rect 42628 6254 42656 6598
rect 42616 6248 42668 6254
rect 42616 6190 42668 6196
rect 42892 6248 42944 6254
rect 42892 6190 42944 6196
rect 42340 6180 42392 6186
rect 42340 6122 42392 6128
rect 42432 6180 42484 6186
rect 42432 6122 42484 6128
rect 42352 5778 42380 6122
rect 42340 5772 42392 5778
rect 42340 5714 42392 5720
rect 42444 5574 42472 6122
rect 42800 6112 42852 6118
rect 42800 6054 42852 6060
rect 42812 5914 42840 6054
rect 42904 5914 42932 6190
rect 42800 5908 42852 5914
rect 42800 5850 42852 5856
rect 42892 5908 42944 5914
rect 42892 5850 42944 5856
rect 42432 5568 42484 5574
rect 42432 5510 42484 5516
rect 42248 5160 42300 5166
rect 42248 5102 42300 5108
rect 41984 4690 42104 4706
rect 41972 4684 42104 4690
rect 42024 4678 42104 4684
rect 41972 4626 42024 4632
rect 43088 4078 43116 7278
rect 43364 7274 43392 9318
rect 43536 7948 43588 7954
rect 43536 7890 43588 7896
rect 43548 7750 43576 7890
rect 43444 7744 43496 7750
rect 43444 7686 43496 7692
rect 43536 7744 43588 7750
rect 43536 7686 43588 7692
rect 43352 7268 43404 7274
rect 43352 7210 43404 7216
rect 43456 6798 43484 7686
rect 43444 6792 43496 6798
rect 43444 6734 43496 6740
rect 43076 4072 43128 4078
rect 43076 4014 43128 4020
rect 41681 3836 41977 3856
rect 41737 3834 41761 3836
rect 41817 3834 41841 3836
rect 41897 3834 41921 3836
rect 41759 3782 41761 3834
rect 41823 3782 41835 3834
rect 41897 3782 41899 3834
rect 41737 3780 41761 3782
rect 41817 3780 41841 3782
rect 41897 3780 41921 3782
rect 41681 3760 41977 3780
rect 41604 3732 41656 3738
rect 41604 3674 41656 3680
rect 43352 3732 43404 3738
rect 43352 3674 43404 3680
rect 42062 3496 42118 3505
rect 42062 3431 42118 3440
rect 41236 3334 41288 3340
rect 41326 3360 41382 3369
rect 41326 3295 41382 3304
rect 41512 3188 41564 3194
rect 41512 3130 41564 3136
rect 40776 3120 40828 3126
rect 40776 3062 40828 3068
rect 39120 3052 39172 3058
rect 39120 2994 39172 3000
rect 38750 2952 38806 2961
rect 38750 2887 38806 2896
rect 40500 2916 40552 2922
rect 40500 2858 40552 2864
rect 37924 2508 37976 2514
rect 37924 2450 37976 2456
rect 38660 2508 38712 2514
rect 38660 2450 38712 2456
rect 40224 2440 40276 2446
rect 40224 2382 40276 2388
rect 39488 2304 39540 2310
rect 39488 2246 39540 2252
rect 37648 2032 37700 2038
rect 37648 1974 37700 1980
rect 36360 1964 36412 1970
rect 36360 1906 36412 1912
rect 36084 1828 36136 1834
rect 36084 1770 36136 1776
rect 36728 1828 36780 1834
rect 36728 1770 36780 1776
rect 36740 800 36768 1770
rect 37660 800 37688 1974
rect 38476 1896 38528 1902
rect 38476 1838 38528 1844
rect 38488 800 38516 1838
rect 39500 1170 39528 2246
rect 39408 1142 39528 1170
rect 39408 800 39436 1142
rect 40236 800 40264 2382
rect 40512 2106 40540 2858
rect 40788 2582 40816 3062
rect 41328 2984 41380 2990
rect 41328 2926 41380 2932
rect 40776 2576 40828 2582
rect 40776 2518 40828 2524
rect 41340 2514 41368 2926
rect 41524 2650 41552 3130
rect 42076 2990 42104 3431
rect 42064 2984 42116 2990
rect 42064 2926 42116 2932
rect 43364 2854 43392 3674
rect 43640 3602 43668 14418
rect 43732 14006 43760 14486
rect 44192 14074 44220 15506
rect 44468 15162 44496 15914
rect 44456 15156 44508 15162
rect 44456 15098 44508 15104
rect 44364 14952 44416 14958
rect 44364 14894 44416 14900
rect 44376 14074 44404 14894
rect 44456 14408 44508 14414
rect 44456 14350 44508 14356
rect 44180 14068 44232 14074
rect 44180 14010 44232 14016
rect 44364 14068 44416 14074
rect 44364 14010 44416 14016
rect 43720 14000 43772 14006
rect 43720 13942 43772 13948
rect 44088 13864 44140 13870
rect 44088 13806 44140 13812
rect 43812 12164 43864 12170
rect 43812 12106 43864 12112
rect 43720 11824 43772 11830
rect 43720 11766 43772 11772
rect 43732 10810 43760 11766
rect 43824 11218 43852 12106
rect 44100 11286 44128 13806
rect 44364 13320 44416 13326
rect 44364 13262 44416 13268
rect 44376 12782 44404 13262
rect 44364 12776 44416 12782
rect 44364 12718 44416 12724
rect 44376 11762 44404 12718
rect 44364 11756 44416 11762
rect 44364 11698 44416 11704
rect 44088 11280 44140 11286
rect 44088 11222 44140 11228
rect 43812 11212 43864 11218
rect 43812 11154 43864 11160
rect 43812 11008 43864 11014
rect 43812 10950 43864 10956
rect 43720 10804 43772 10810
rect 43720 10746 43772 10752
rect 43732 10198 43760 10746
rect 43720 10192 43772 10198
rect 43720 10134 43772 10140
rect 43720 5160 43772 5166
rect 43720 5102 43772 5108
rect 43732 4826 43760 5102
rect 43720 4820 43772 4826
rect 43720 4762 43772 4768
rect 43628 3596 43680 3602
rect 43628 3538 43680 3544
rect 43824 3466 43852 10950
rect 44468 10146 44496 14350
rect 44560 12374 44588 15982
rect 44744 14890 44772 15982
rect 45020 14958 45048 17274
rect 46204 17060 46256 17066
rect 46204 17002 46256 17008
rect 45928 16652 45980 16658
rect 45928 16594 45980 16600
rect 45192 15904 45244 15910
rect 45192 15846 45244 15852
rect 45204 15638 45232 15846
rect 45192 15632 45244 15638
rect 45192 15574 45244 15580
rect 45284 15564 45336 15570
rect 45284 15506 45336 15512
rect 45008 14952 45060 14958
rect 45008 14894 45060 14900
rect 44732 14884 44784 14890
rect 44732 14826 44784 14832
rect 44732 13864 44784 13870
rect 44732 13806 44784 13812
rect 44916 13864 44968 13870
rect 44916 13806 44968 13812
rect 44744 13326 44772 13806
rect 44732 13320 44784 13326
rect 44732 13262 44784 13268
rect 44548 12368 44600 12374
rect 44548 12310 44600 12316
rect 44744 12238 44772 13262
rect 44732 12232 44784 12238
rect 44732 12174 44784 12180
rect 44824 11144 44876 11150
rect 44824 11086 44876 11092
rect 44836 10606 44864 11086
rect 44824 10600 44876 10606
rect 44824 10542 44876 10548
rect 44928 10266 44956 13806
rect 45296 13462 45324 15506
rect 45940 14482 45968 16594
rect 46112 16584 46164 16590
rect 46112 16526 46164 16532
rect 46124 15638 46152 16526
rect 46216 16046 46244 17002
rect 46952 16794 46980 18835
rect 48884 17134 48912 18835
rect 50816 17134 50844 18835
rect 51862 17436 52158 17456
rect 51918 17434 51942 17436
rect 51998 17434 52022 17436
rect 52078 17434 52102 17436
rect 51940 17382 51942 17434
rect 52004 17382 52016 17434
rect 52078 17382 52080 17434
rect 51918 17380 51942 17382
rect 51998 17380 52022 17382
rect 52078 17380 52102 17382
rect 51862 17360 52158 17380
rect 48872 17128 48924 17134
rect 48872 17070 48924 17076
rect 50804 17128 50856 17134
rect 50804 17070 50856 17076
rect 48504 16992 48556 16998
rect 48504 16934 48556 16940
rect 46940 16788 46992 16794
rect 46940 16730 46992 16736
rect 46664 16108 46716 16114
rect 46664 16050 46716 16056
rect 46204 16040 46256 16046
rect 46204 15982 46256 15988
rect 46112 15632 46164 15638
rect 46112 15574 46164 15580
rect 46676 14958 46704 16050
rect 46952 16046 46980 16730
rect 48044 16652 48096 16658
rect 48044 16594 48096 16600
rect 48056 16046 48084 16594
rect 46940 16040 46992 16046
rect 46940 15982 46992 15988
rect 48044 16040 48096 16046
rect 48044 15982 48096 15988
rect 48320 16040 48372 16046
rect 48320 15982 48372 15988
rect 46940 15564 46992 15570
rect 46940 15506 46992 15512
rect 46664 14952 46716 14958
rect 46664 14894 46716 14900
rect 46296 14816 46348 14822
rect 46296 14758 46348 14764
rect 45928 14476 45980 14482
rect 45928 14418 45980 14424
rect 46112 14476 46164 14482
rect 46112 14418 46164 14424
rect 45468 14272 45520 14278
rect 45468 14214 45520 14220
rect 45284 13456 45336 13462
rect 45284 13398 45336 13404
rect 45100 12844 45152 12850
rect 45100 12786 45152 12792
rect 45112 10674 45140 12786
rect 45376 12776 45428 12782
rect 45376 12718 45428 12724
rect 45192 12300 45244 12306
rect 45192 12242 45244 12248
rect 45204 11898 45232 12242
rect 45192 11892 45244 11898
rect 45192 11834 45244 11840
rect 45284 11824 45336 11830
rect 45284 11766 45336 11772
rect 45190 11656 45246 11665
rect 45190 11591 45192 11600
rect 45244 11591 45246 11600
rect 45192 11562 45244 11568
rect 45296 11234 45324 11766
rect 45204 11206 45324 11234
rect 45204 11150 45232 11206
rect 45192 11144 45244 11150
rect 45192 11086 45244 11092
rect 45100 10668 45152 10674
rect 45100 10610 45152 10616
rect 44916 10260 44968 10266
rect 44916 10202 44968 10208
rect 44468 10118 44772 10146
rect 44468 9738 44496 10118
rect 44640 10056 44692 10062
rect 44640 9998 44692 10004
rect 44376 9722 44496 9738
rect 44364 9716 44496 9722
rect 44416 9710 44496 9716
rect 44364 9658 44416 9664
rect 43904 9580 43956 9586
rect 43904 9522 43956 9528
rect 43916 6866 43944 9522
rect 44364 9512 44416 9518
rect 44364 9454 44416 9460
rect 44088 9444 44140 9450
rect 44088 9386 44140 9392
rect 44100 9330 44128 9386
rect 44100 9302 44220 9330
rect 44192 9081 44220 9302
rect 44178 9072 44234 9081
rect 44178 9007 44234 9016
rect 44272 9036 44324 9042
rect 44272 8978 44324 8984
rect 43996 8968 44048 8974
rect 43996 8910 44048 8916
rect 44008 8022 44036 8910
rect 44180 8424 44232 8430
rect 44180 8366 44232 8372
rect 44192 8265 44220 8366
rect 44178 8256 44234 8265
rect 44178 8191 44234 8200
rect 43996 8016 44048 8022
rect 43996 7958 44048 7964
rect 44008 7342 44036 7958
rect 44088 7948 44140 7954
rect 44088 7890 44140 7896
rect 44100 7546 44128 7890
rect 44088 7540 44140 7546
rect 44088 7482 44140 7488
rect 44284 7410 44312 8978
rect 44376 8430 44404 9454
rect 44456 8832 44508 8838
rect 44456 8774 44508 8780
rect 44468 8430 44496 8774
rect 44652 8634 44680 9998
rect 44744 9364 44772 10118
rect 44928 9722 44956 10202
rect 45100 10124 45152 10130
rect 45204 10112 45232 11086
rect 45152 10084 45232 10112
rect 45100 10066 45152 10072
rect 44916 9716 44968 9722
rect 44916 9658 44968 9664
rect 45192 9716 45244 9722
rect 45192 9658 45244 9664
rect 45008 9376 45060 9382
rect 44744 9336 45008 9364
rect 45008 9318 45060 9324
rect 44916 9036 44968 9042
rect 44916 8978 44968 8984
rect 44824 8900 44876 8906
rect 44824 8842 44876 8848
rect 44640 8628 44692 8634
rect 44640 8570 44692 8576
rect 44836 8430 44864 8842
rect 44364 8424 44416 8430
rect 44364 8366 44416 8372
rect 44456 8424 44508 8430
rect 44456 8366 44508 8372
rect 44824 8424 44876 8430
rect 44824 8366 44876 8372
rect 44824 8288 44876 8294
rect 44824 8230 44876 8236
rect 44456 7948 44508 7954
rect 44456 7890 44508 7896
rect 44272 7404 44324 7410
rect 44272 7346 44324 7352
rect 43996 7336 44048 7342
rect 43996 7278 44048 7284
rect 44284 6866 44312 7346
rect 44468 7313 44496 7890
rect 44732 7880 44784 7886
rect 44732 7822 44784 7828
rect 44744 7410 44772 7822
rect 44732 7404 44784 7410
rect 44732 7346 44784 7352
rect 44454 7304 44510 7313
rect 44454 7239 44510 7248
rect 43904 6860 43956 6866
rect 43904 6802 43956 6808
rect 44272 6860 44324 6866
rect 44272 6802 44324 6808
rect 44364 6792 44416 6798
rect 44362 6760 44364 6769
rect 44416 6760 44418 6769
rect 44362 6695 44418 6704
rect 44468 5778 44496 7239
rect 44744 7206 44772 7346
rect 44732 7200 44784 7206
rect 44732 7142 44784 7148
rect 44836 6304 44864 8230
rect 44928 8090 44956 8978
rect 45204 8838 45232 9658
rect 45388 9081 45416 12718
rect 45374 9072 45430 9081
rect 45480 9042 45508 14214
rect 45652 13864 45704 13870
rect 45652 13806 45704 13812
rect 45664 13326 45692 13806
rect 45744 13388 45796 13394
rect 45744 13330 45796 13336
rect 45652 13320 45704 13326
rect 45652 13262 45704 13268
rect 45560 12300 45612 12306
rect 45560 12242 45612 12248
rect 45572 9586 45600 12242
rect 45560 9580 45612 9586
rect 45612 9540 45692 9568
rect 45560 9522 45612 9528
rect 45664 9110 45692 9540
rect 45652 9104 45704 9110
rect 45652 9046 45704 9052
rect 45374 9007 45430 9016
rect 45468 9036 45520 9042
rect 45468 8978 45520 8984
rect 45756 8974 45784 13330
rect 45836 13320 45888 13326
rect 45836 13262 45888 13268
rect 45848 12306 45876 13262
rect 45940 13190 45968 14418
rect 46124 14074 46152 14418
rect 46112 14068 46164 14074
rect 46112 14010 46164 14016
rect 46308 13802 46336 14758
rect 46676 14550 46704 14894
rect 46664 14544 46716 14550
rect 46664 14486 46716 14492
rect 46572 14408 46624 14414
rect 46572 14350 46624 14356
rect 46584 14074 46612 14350
rect 46572 14068 46624 14074
rect 46572 14010 46624 14016
rect 46388 13864 46440 13870
rect 46388 13806 46440 13812
rect 46296 13796 46348 13802
rect 46296 13738 46348 13744
rect 46204 13728 46256 13734
rect 46204 13670 46256 13676
rect 46112 13388 46164 13394
rect 46112 13330 46164 13336
rect 45928 13184 45980 13190
rect 45928 13126 45980 13132
rect 46124 12986 46152 13330
rect 46112 12980 46164 12986
rect 46112 12922 46164 12928
rect 46216 12458 46244 13670
rect 46400 12986 46428 13806
rect 46952 13258 46980 15506
rect 47032 15020 47084 15026
rect 47032 14962 47084 14968
rect 47044 13870 47072 14962
rect 47216 14612 47268 14618
rect 47216 14554 47268 14560
rect 47032 13864 47084 13870
rect 47032 13806 47084 13812
rect 46480 13252 46532 13258
rect 46480 13194 46532 13200
rect 46940 13252 46992 13258
rect 46940 13194 46992 13200
rect 46388 12980 46440 12986
rect 46388 12922 46440 12928
rect 46216 12430 46336 12458
rect 45836 12300 45888 12306
rect 45836 12242 45888 12248
rect 46204 12164 46256 12170
rect 46204 12106 46256 12112
rect 46216 11694 46244 12106
rect 46308 12050 46336 12430
rect 46308 12022 46428 12050
rect 46294 11928 46350 11937
rect 46294 11863 46350 11872
rect 46308 11762 46336 11863
rect 46296 11756 46348 11762
rect 46296 11698 46348 11704
rect 46204 11688 46256 11694
rect 46204 11630 46256 11636
rect 46112 11144 46164 11150
rect 46112 11086 46164 11092
rect 46124 10674 46152 11086
rect 46112 10668 46164 10674
rect 46112 10610 46164 10616
rect 45928 10600 45980 10606
rect 45928 10542 45980 10548
rect 45744 8968 45796 8974
rect 45744 8910 45796 8916
rect 45192 8832 45244 8838
rect 45192 8774 45244 8780
rect 45836 8832 45888 8838
rect 45836 8774 45888 8780
rect 44916 8084 44968 8090
rect 44916 8026 44968 8032
rect 44928 6798 44956 8026
rect 45204 7342 45232 8774
rect 45848 8430 45876 8774
rect 45836 8424 45888 8430
rect 45296 8350 45600 8378
rect 45836 8366 45888 8372
rect 45296 7886 45324 8350
rect 45572 8294 45600 8350
rect 45560 8288 45612 8294
rect 45560 8230 45612 8236
rect 45284 7880 45336 7886
rect 45284 7822 45336 7828
rect 45560 7880 45612 7886
rect 45744 7880 45796 7886
rect 45560 7822 45612 7828
rect 45742 7848 45744 7857
rect 45796 7848 45798 7857
rect 45192 7336 45244 7342
rect 45192 7278 45244 7284
rect 45572 7002 45600 7822
rect 45742 7783 45798 7792
rect 45560 6996 45612 7002
rect 45560 6938 45612 6944
rect 45652 6860 45704 6866
rect 45652 6802 45704 6808
rect 44916 6792 44968 6798
rect 44916 6734 44968 6740
rect 44916 6316 44968 6322
rect 44836 6276 44916 6304
rect 44916 6258 44968 6264
rect 44640 6248 44692 6254
rect 44640 6190 44692 6196
rect 44652 5846 44680 6190
rect 44640 5840 44692 5846
rect 44640 5782 44692 5788
rect 44088 5772 44140 5778
rect 44088 5714 44140 5720
rect 44456 5772 44508 5778
rect 44456 5714 44508 5720
rect 44100 5658 44128 5714
rect 44100 5630 44220 5658
rect 44192 5098 44220 5630
rect 44180 5092 44232 5098
rect 44180 5034 44232 5040
rect 44928 4078 44956 6258
rect 45560 6112 45612 6118
rect 45560 6054 45612 6060
rect 45190 5808 45246 5817
rect 45190 5743 45246 5752
rect 45204 5710 45232 5743
rect 45192 5704 45244 5710
rect 45192 5646 45244 5652
rect 45468 5704 45520 5710
rect 45468 5646 45520 5652
rect 45480 5234 45508 5646
rect 45468 5228 45520 5234
rect 45468 5170 45520 5176
rect 45468 4684 45520 4690
rect 45468 4626 45520 4632
rect 45480 4078 45508 4626
rect 45572 4146 45600 6054
rect 45664 5817 45692 6802
rect 45650 5808 45706 5817
rect 45650 5743 45652 5752
rect 45704 5743 45706 5752
rect 45652 5714 45704 5720
rect 45652 5636 45704 5642
rect 45652 5578 45704 5584
rect 45560 4140 45612 4146
rect 45560 4082 45612 4088
rect 44916 4072 44968 4078
rect 44916 4014 44968 4020
rect 45468 4072 45520 4078
rect 45468 4014 45520 4020
rect 45664 3942 45692 5578
rect 45756 4826 45784 7783
rect 45940 6497 45968 10542
rect 46400 10470 46428 12022
rect 46388 10464 46440 10470
rect 46388 10406 46440 10412
rect 46112 10124 46164 10130
rect 46112 10066 46164 10072
rect 46124 9586 46152 10066
rect 46112 9580 46164 9586
rect 46112 9522 46164 9528
rect 46400 9518 46428 10406
rect 46388 9512 46440 9518
rect 46388 9454 46440 9460
rect 46492 9450 46520 13194
rect 46664 13184 46716 13190
rect 46664 13126 46716 13132
rect 46572 12232 46624 12238
rect 46572 12174 46624 12180
rect 46584 11014 46612 12174
rect 46676 11830 46704 13126
rect 47044 12918 47072 13806
rect 47228 13802 47256 14554
rect 48056 14482 48084 15982
rect 48332 15638 48360 15982
rect 48516 15706 48544 16934
rect 48884 16266 48912 17070
rect 49976 16992 50028 16998
rect 49976 16934 50028 16940
rect 49700 16584 49752 16590
rect 49700 16526 49752 16532
rect 48884 16250 49004 16266
rect 48884 16244 49016 16250
rect 48884 16238 48964 16244
rect 48964 16186 49016 16192
rect 48504 15700 48556 15706
rect 48504 15642 48556 15648
rect 49712 15638 49740 16526
rect 49988 15706 50016 16934
rect 50816 16794 50844 17070
rect 50804 16788 50856 16794
rect 50804 16730 50856 16736
rect 51862 16348 52158 16368
rect 51918 16346 51942 16348
rect 51998 16346 52022 16348
rect 52078 16346 52102 16348
rect 51940 16294 51942 16346
rect 52004 16294 52016 16346
rect 52078 16294 52080 16346
rect 51918 16292 51942 16294
rect 51998 16292 52022 16294
rect 52078 16292 52102 16294
rect 51862 16272 52158 16292
rect 49976 15700 50028 15706
rect 49976 15642 50028 15648
rect 52656 15638 52684 18835
rect 48320 15632 48372 15638
rect 48320 15574 48372 15580
rect 49700 15632 49752 15638
rect 49700 15574 49752 15580
rect 51632 15632 51684 15638
rect 51632 15574 51684 15580
rect 52644 15632 52696 15638
rect 52644 15574 52696 15580
rect 49240 15564 49292 15570
rect 49240 15506 49292 15512
rect 49608 15564 49660 15570
rect 49608 15506 49660 15512
rect 48044 14476 48096 14482
rect 48044 14418 48096 14424
rect 47400 13932 47452 13938
rect 47400 13874 47452 13880
rect 48228 13932 48280 13938
rect 48228 13874 48280 13880
rect 47216 13796 47268 13802
rect 47216 13738 47268 13744
rect 47124 13388 47176 13394
rect 47124 13330 47176 13336
rect 47032 12912 47084 12918
rect 47032 12854 47084 12860
rect 47032 12776 47084 12782
rect 47032 12718 47084 12724
rect 46664 11824 46716 11830
rect 46664 11766 46716 11772
rect 46572 11008 46624 11014
rect 46572 10950 46624 10956
rect 46940 11008 46992 11014
rect 46940 10950 46992 10956
rect 46952 10606 46980 10950
rect 46940 10600 46992 10606
rect 46940 10542 46992 10548
rect 46112 9444 46164 9450
rect 46112 9386 46164 9392
rect 46480 9444 46532 9450
rect 46480 9386 46532 9392
rect 46848 9444 46900 9450
rect 46848 9386 46900 9392
rect 46124 8362 46152 9386
rect 46204 9376 46256 9382
rect 46204 9318 46256 9324
rect 46216 8548 46244 9318
rect 46296 8560 46348 8566
rect 46216 8520 46296 8548
rect 46112 8356 46164 8362
rect 46112 8298 46164 8304
rect 46020 8288 46072 8294
rect 46020 8230 46072 8236
rect 46032 6644 46060 8230
rect 46216 8090 46244 8520
rect 46296 8502 46348 8508
rect 46860 8430 46888 9386
rect 47044 9058 47072 12718
rect 47136 12374 47164 13330
rect 47228 12850 47256 13738
rect 47412 13326 47440 13874
rect 48136 13728 48188 13734
rect 48136 13670 48188 13676
rect 48148 13394 48176 13670
rect 47584 13388 47636 13394
rect 47584 13330 47636 13336
rect 48136 13388 48188 13394
rect 48136 13330 48188 13336
rect 47400 13320 47452 13326
rect 47400 13262 47452 13268
rect 47216 12844 47268 12850
rect 47216 12786 47268 12792
rect 47124 12368 47176 12374
rect 47124 12310 47176 12316
rect 47492 11348 47544 11354
rect 47492 11290 47544 11296
rect 47504 11150 47532 11290
rect 47492 11144 47544 11150
rect 47492 11086 47544 11092
rect 47216 10600 47268 10606
rect 47216 10542 47268 10548
rect 47228 10198 47256 10542
rect 47492 10260 47544 10266
rect 47492 10202 47544 10208
rect 47216 10192 47268 10198
rect 47216 10134 47268 10140
rect 47044 9030 47164 9058
rect 46940 8968 46992 8974
rect 46940 8910 46992 8916
rect 46952 8498 46980 8910
rect 46940 8492 46992 8498
rect 46940 8434 46992 8440
rect 46296 8424 46348 8430
rect 46296 8366 46348 8372
rect 46848 8424 46900 8430
rect 46848 8366 46900 8372
rect 46112 8084 46164 8090
rect 46112 8026 46164 8032
rect 46204 8084 46256 8090
rect 46204 8026 46256 8032
rect 46124 7954 46152 8026
rect 46112 7948 46164 7954
rect 46112 7890 46164 7896
rect 46216 7342 46244 8026
rect 46204 7336 46256 7342
rect 46204 7278 46256 7284
rect 46112 7268 46164 7274
rect 46112 7210 46164 7216
rect 46124 6798 46152 7210
rect 46112 6792 46164 6798
rect 46112 6734 46164 6740
rect 46032 6616 46152 6644
rect 45926 6488 45982 6497
rect 45926 6423 45982 6432
rect 46124 5166 46152 6616
rect 46308 6304 46336 8366
rect 46388 8288 46440 8294
rect 46388 8230 46440 8236
rect 46400 7410 46428 8230
rect 47136 7698 47164 9030
rect 47228 7750 47256 10134
rect 47504 9518 47532 10202
rect 47492 9512 47544 9518
rect 47492 9454 47544 9460
rect 47306 8800 47362 8809
rect 47306 8735 47362 8744
rect 47044 7670 47164 7698
rect 47216 7744 47268 7750
rect 47216 7686 47268 7692
rect 46388 7404 46440 7410
rect 46388 7346 46440 7352
rect 47044 6866 47072 7670
rect 47320 7449 47348 8735
rect 47492 7948 47544 7954
rect 47492 7890 47544 7896
rect 47504 7478 47532 7890
rect 47492 7472 47544 7478
rect 47306 7440 47362 7449
rect 47216 7404 47268 7410
rect 47492 7414 47544 7420
rect 47306 7375 47362 7384
rect 47216 7346 47268 7352
rect 47228 7206 47256 7346
rect 47216 7200 47268 7206
rect 47216 7142 47268 7148
rect 47306 6896 47362 6905
rect 46756 6860 46808 6866
rect 46756 6802 46808 6808
rect 47032 6860 47084 6866
rect 47306 6831 47362 6840
rect 47032 6802 47084 6808
rect 46572 6792 46624 6798
rect 46572 6734 46624 6740
rect 46216 6276 46336 6304
rect 46216 5166 46244 6276
rect 46584 6202 46612 6734
rect 46308 6186 46612 6202
rect 46296 6180 46612 6186
rect 46348 6174 46612 6180
rect 46296 6122 46348 6128
rect 46388 5704 46440 5710
rect 46388 5646 46440 5652
rect 46400 5234 46428 5646
rect 46388 5228 46440 5234
rect 46388 5170 46440 5176
rect 46112 5160 46164 5166
rect 46112 5102 46164 5108
rect 46204 5160 46256 5166
rect 46204 5102 46256 5108
rect 45744 4820 45796 4826
rect 45744 4762 45796 4768
rect 45756 4214 45784 4762
rect 45744 4208 45796 4214
rect 45744 4150 45796 4156
rect 45652 3936 45704 3942
rect 45652 3878 45704 3884
rect 44088 3596 44140 3602
rect 44088 3538 44140 3544
rect 43812 3460 43864 3466
rect 43812 3402 43864 3408
rect 44100 2854 44128 3538
rect 46124 3534 46152 5102
rect 46584 4690 46612 6174
rect 46768 6118 46796 6802
rect 46848 6724 46900 6730
rect 46848 6666 46900 6672
rect 46756 6112 46808 6118
rect 46756 6054 46808 6060
rect 46754 5536 46810 5545
rect 46754 5471 46810 5480
rect 46768 5137 46796 5471
rect 46754 5128 46810 5137
rect 46754 5063 46810 5072
rect 46572 4684 46624 4690
rect 46572 4626 46624 4632
rect 46860 4282 46888 6666
rect 47044 6662 47072 6802
rect 47320 6798 47348 6831
rect 47308 6792 47360 6798
rect 47308 6734 47360 6740
rect 47032 6656 47084 6662
rect 47032 6598 47084 6604
rect 47216 5908 47268 5914
rect 47216 5850 47268 5856
rect 47228 5642 47256 5850
rect 47216 5636 47268 5642
rect 47216 5578 47268 5584
rect 47490 5264 47546 5273
rect 47596 5250 47624 13330
rect 48240 13326 48268 13874
rect 49252 13462 49280 15506
rect 49620 15162 49648 15506
rect 51540 15496 51592 15502
rect 51540 15438 51592 15444
rect 49608 15156 49660 15162
rect 49608 15098 49660 15104
rect 50252 15020 50304 15026
rect 50252 14962 50304 14968
rect 50264 14482 50292 14962
rect 50252 14476 50304 14482
rect 50252 14418 50304 14424
rect 51552 13938 51580 15438
rect 51644 14618 51672 15574
rect 53288 15564 53340 15570
rect 53288 15506 53340 15512
rect 52920 15496 52972 15502
rect 52920 15438 52972 15444
rect 51862 15260 52158 15280
rect 51918 15258 51942 15260
rect 51998 15258 52022 15260
rect 52078 15258 52102 15260
rect 51940 15206 51942 15258
rect 52004 15206 52016 15258
rect 52078 15206 52080 15258
rect 51918 15204 51942 15206
rect 51998 15204 52022 15206
rect 52078 15204 52102 15206
rect 51862 15184 52158 15204
rect 51632 14612 51684 14618
rect 51632 14554 51684 14560
rect 52932 14550 52960 15438
rect 53300 15366 53328 15506
rect 54588 15366 54616 18835
rect 55312 16652 55364 16658
rect 55312 16594 55364 16600
rect 55588 16652 55640 16658
rect 55588 16594 55640 16600
rect 55128 15972 55180 15978
rect 55128 15914 55180 15920
rect 55140 15434 55168 15914
rect 54668 15428 54720 15434
rect 54668 15370 54720 15376
rect 55128 15428 55180 15434
rect 55128 15370 55180 15376
rect 53288 15360 53340 15366
rect 53288 15302 53340 15308
rect 54576 15360 54628 15366
rect 54576 15302 54628 15308
rect 53300 15162 53328 15302
rect 53288 15156 53340 15162
rect 53288 15098 53340 15104
rect 53472 14952 53524 14958
rect 53472 14894 53524 14900
rect 53484 14550 53512 14894
rect 52920 14544 52972 14550
rect 52920 14486 52972 14492
rect 53472 14544 53524 14550
rect 53472 14486 53524 14492
rect 53012 14476 53064 14482
rect 53012 14418 53064 14424
rect 52184 14408 52236 14414
rect 52184 14350 52236 14356
rect 51862 14172 52158 14192
rect 51918 14170 51942 14172
rect 51998 14170 52022 14172
rect 52078 14170 52102 14172
rect 51940 14118 51942 14170
rect 52004 14118 52016 14170
rect 52078 14118 52080 14170
rect 51918 14116 51942 14118
rect 51998 14116 52022 14118
rect 52078 14116 52102 14118
rect 51862 14096 52158 14116
rect 52196 14074 52224 14350
rect 52736 14272 52788 14278
rect 52736 14214 52788 14220
rect 52748 14074 52776 14214
rect 52184 14068 52236 14074
rect 52184 14010 52236 14016
rect 52736 14068 52788 14074
rect 52736 14010 52788 14016
rect 51540 13932 51592 13938
rect 51540 13874 51592 13880
rect 52552 13864 52604 13870
rect 52552 13806 52604 13812
rect 50068 13728 50120 13734
rect 50068 13670 50120 13676
rect 49240 13456 49292 13462
rect 49240 13398 49292 13404
rect 49608 13388 49660 13394
rect 49608 13330 49660 13336
rect 49976 13388 50028 13394
rect 49976 13330 50028 13336
rect 48228 13320 48280 13326
rect 48228 13262 48280 13268
rect 49620 12986 49648 13330
rect 49608 12980 49660 12986
rect 49608 12922 49660 12928
rect 48228 12912 48280 12918
rect 48228 12854 48280 12860
rect 48136 12776 48188 12782
rect 48136 12718 48188 12724
rect 48044 12708 48096 12714
rect 48044 12650 48096 12656
rect 48056 11286 48084 12650
rect 48044 11280 48096 11286
rect 48044 11222 48096 11228
rect 48148 10577 48176 12718
rect 48240 12306 48268 12854
rect 48228 12300 48280 12306
rect 48228 12242 48280 12248
rect 49700 11892 49752 11898
rect 49700 11834 49752 11840
rect 49240 11824 49292 11830
rect 49240 11766 49292 11772
rect 48780 11688 48832 11694
rect 48686 11656 48742 11665
rect 48780 11630 48832 11636
rect 48686 11591 48688 11600
rect 48740 11591 48742 11600
rect 48688 11562 48740 11568
rect 48412 11008 48464 11014
rect 48412 10950 48464 10956
rect 48134 10568 48190 10577
rect 48424 10538 48452 10950
rect 48134 10503 48190 10512
rect 48412 10532 48464 10538
rect 48148 9722 48176 10503
rect 48412 10474 48464 10480
rect 48136 9716 48188 9722
rect 48136 9658 48188 9664
rect 48596 9716 48648 9722
rect 48596 9658 48648 9664
rect 48504 9648 48556 9654
rect 48504 9590 48556 9596
rect 47768 9512 47820 9518
rect 47768 9454 47820 9460
rect 47780 8888 47808 9454
rect 48516 9081 48544 9590
rect 47950 9072 48006 9081
rect 47950 9007 47952 9016
rect 48004 9007 48006 9016
rect 48502 9072 48558 9081
rect 48502 9007 48558 9016
rect 47952 8978 48004 8984
rect 47860 8900 47912 8906
rect 47780 8860 47860 8888
rect 47780 8090 47808 8860
rect 47860 8842 47912 8848
rect 48410 8800 48466 8809
rect 48410 8735 48466 8744
rect 47964 8634 48176 8650
rect 47964 8628 48188 8634
rect 47964 8622 48136 8628
rect 47964 8362 47992 8622
rect 48136 8570 48188 8576
rect 48424 8498 48452 8735
rect 48412 8492 48464 8498
rect 48412 8434 48464 8440
rect 47952 8356 48004 8362
rect 47952 8298 48004 8304
rect 47768 8084 47820 8090
rect 47768 8026 47820 8032
rect 48228 7200 48280 7206
rect 48228 7142 48280 7148
rect 47964 6718 48176 6746
rect 47964 6662 47992 6718
rect 47952 6656 48004 6662
rect 47952 6598 48004 6604
rect 48044 6656 48096 6662
rect 48044 6598 48096 6604
rect 48056 5710 48084 6598
rect 48148 5710 48176 6718
rect 48044 5704 48096 5710
rect 48044 5646 48096 5652
rect 48136 5704 48188 5710
rect 48136 5646 48188 5652
rect 47676 5636 47728 5642
rect 47676 5578 47728 5584
rect 47688 5302 47716 5578
rect 47546 5222 47624 5250
rect 47676 5296 47728 5302
rect 47676 5238 47728 5244
rect 47490 5199 47546 5208
rect 46938 5128 46994 5137
rect 46938 5063 46994 5072
rect 46952 4486 46980 5063
rect 46940 4480 46992 4486
rect 46940 4422 46992 4428
rect 46848 4276 46900 4282
rect 46848 4218 46900 4224
rect 47596 4078 47624 5222
rect 47952 5092 48004 5098
rect 47952 5034 48004 5040
rect 47964 4758 47992 5034
rect 47952 4752 48004 4758
rect 47952 4694 48004 4700
rect 47584 4072 47636 4078
rect 47584 4014 47636 4020
rect 46572 4004 46624 4010
rect 46572 3946 46624 3952
rect 46584 3602 46612 3946
rect 46572 3596 46624 3602
rect 46572 3538 46624 3544
rect 46112 3528 46164 3534
rect 46112 3470 46164 3476
rect 47032 3188 47084 3194
rect 47032 3130 47084 3136
rect 47044 2990 47072 3130
rect 47596 2990 47624 4014
rect 48240 4010 48268 7142
rect 48318 6896 48374 6905
rect 48318 6831 48374 6840
rect 48332 6458 48360 6831
rect 48320 6452 48372 6458
rect 48320 6394 48372 6400
rect 48228 4004 48280 4010
rect 48228 3946 48280 3952
rect 45192 2984 45244 2990
rect 45192 2926 45244 2932
rect 47032 2984 47084 2990
rect 47032 2926 47084 2932
rect 47584 2984 47636 2990
rect 47584 2926 47636 2932
rect 44640 2916 44692 2922
rect 44640 2858 44692 2864
rect 43352 2848 43404 2854
rect 43352 2790 43404 2796
rect 44088 2848 44140 2854
rect 44088 2790 44140 2796
rect 41681 2748 41977 2768
rect 41737 2746 41761 2748
rect 41817 2746 41841 2748
rect 41897 2746 41921 2748
rect 41759 2694 41761 2746
rect 41823 2694 41835 2746
rect 41897 2694 41899 2746
rect 41737 2692 41761 2694
rect 41817 2692 41841 2694
rect 41897 2692 41921 2694
rect 41681 2672 41977 2692
rect 44652 2650 44680 2858
rect 45204 2650 45232 2926
rect 48504 2848 48556 2854
rect 48504 2790 48556 2796
rect 41512 2644 41564 2650
rect 41512 2586 41564 2592
rect 44640 2644 44692 2650
rect 44640 2586 44692 2592
rect 45192 2644 45244 2650
rect 45192 2586 45244 2592
rect 48516 2514 48544 2790
rect 48608 2650 48636 9658
rect 48688 9648 48740 9654
rect 48688 9590 48740 9596
rect 48700 8974 48728 9590
rect 48688 8968 48740 8974
rect 48688 8910 48740 8916
rect 48688 6792 48740 6798
rect 48688 6734 48740 6740
rect 48700 6254 48728 6734
rect 48688 6248 48740 6254
rect 48688 6190 48740 6196
rect 48700 3233 48728 6190
rect 48792 4622 48820 11630
rect 49252 11218 49280 11766
rect 49712 11694 49740 11834
rect 49700 11688 49752 11694
rect 49700 11630 49752 11636
rect 49056 11212 49108 11218
rect 49056 11154 49108 11160
rect 49240 11212 49292 11218
rect 49240 11154 49292 11160
rect 49068 10810 49096 11154
rect 49056 10804 49108 10810
rect 49056 10746 49108 10752
rect 48964 10600 49016 10606
rect 48964 10542 49016 10548
rect 48976 10198 49004 10542
rect 48964 10192 49016 10198
rect 48964 10134 49016 10140
rect 49068 9722 49096 10746
rect 49332 10532 49384 10538
rect 49332 10474 49384 10480
rect 49344 10266 49372 10474
rect 49332 10260 49384 10266
rect 49332 10202 49384 10208
rect 49516 10124 49568 10130
rect 49516 10066 49568 10072
rect 49056 9716 49108 9722
rect 49056 9658 49108 9664
rect 48872 6248 48924 6254
rect 48872 6190 48924 6196
rect 48884 5914 48912 6190
rect 48872 5908 48924 5914
rect 48872 5850 48924 5856
rect 49068 4690 49096 9658
rect 49240 9512 49292 9518
rect 49240 9454 49292 9460
rect 49252 8838 49280 9454
rect 49424 9376 49476 9382
rect 49424 9318 49476 9324
rect 49436 8838 49464 9318
rect 49240 8832 49292 8838
rect 49240 8774 49292 8780
rect 49424 8832 49476 8838
rect 49424 8774 49476 8780
rect 49528 6798 49556 10066
rect 49712 10062 49740 11630
rect 49988 11558 50016 13330
rect 50080 13326 50108 13670
rect 51092 13394 51212 13410
rect 51092 13388 51224 13394
rect 51092 13382 51172 13388
rect 50068 13320 50120 13326
rect 50068 13262 50120 13268
rect 50620 13320 50672 13326
rect 50620 13262 50672 13268
rect 50252 12776 50304 12782
rect 50252 12718 50304 12724
rect 50068 12708 50120 12714
rect 50068 12650 50120 12656
rect 49976 11552 50028 11558
rect 49976 11494 50028 11500
rect 50080 10810 50108 12650
rect 50264 12102 50292 12718
rect 50528 12368 50580 12374
rect 50528 12310 50580 12316
rect 50252 12096 50304 12102
rect 50252 12038 50304 12044
rect 50068 10804 50120 10810
rect 50068 10746 50120 10752
rect 50080 10130 50108 10746
rect 50068 10124 50120 10130
rect 50068 10066 50120 10072
rect 49700 10056 49752 10062
rect 49700 9998 49752 10004
rect 50264 9926 50292 12038
rect 50540 11694 50568 12310
rect 50528 11688 50580 11694
rect 50528 11630 50580 11636
rect 50632 11626 50660 13262
rect 51092 12782 51120 13382
rect 51172 13330 51224 13336
rect 51632 13320 51684 13326
rect 51632 13262 51684 13268
rect 51644 12782 51672 13262
rect 51862 13084 52158 13104
rect 51918 13082 51942 13084
rect 51998 13082 52022 13084
rect 52078 13082 52102 13084
rect 51940 13030 51942 13082
rect 52004 13030 52016 13082
rect 52078 13030 52080 13082
rect 51918 13028 51942 13030
rect 51998 13028 52022 13030
rect 52078 13028 52102 13030
rect 51862 13008 52158 13028
rect 51080 12776 51132 12782
rect 51080 12718 51132 12724
rect 51632 12776 51684 12782
rect 51632 12718 51684 12724
rect 50896 12708 50948 12714
rect 50896 12650 50948 12656
rect 50908 12306 50936 12650
rect 50896 12300 50948 12306
rect 50896 12242 50948 12248
rect 50620 11620 50672 11626
rect 50620 11562 50672 11568
rect 50528 11552 50580 11558
rect 50528 11494 50580 11500
rect 50252 9920 50304 9926
rect 50252 9862 50304 9868
rect 49792 9512 49844 9518
rect 49792 9454 49844 9460
rect 50436 9512 50488 9518
rect 50436 9454 50488 9460
rect 49608 9036 49660 9042
rect 49608 8978 49660 8984
rect 49620 8906 49648 8978
rect 49608 8900 49660 8906
rect 49608 8842 49660 8848
rect 49620 8294 49648 8842
rect 49608 8288 49660 8294
rect 49608 8230 49660 8236
rect 49804 7886 49832 9454
rect 50448 9042 50476 9454
rect 50436 9036 50488 9042
rect 50436 8978 50488 8984
rect 50250 8664 50306 8673
rect 50250 8599 50306 8608
rect 50344 8628 50396 8634
rect 50264 8430 50292 8599
rect 50344 8570 50396 8576
rect 50436 8628 50488 8634
rect 50436 8570 50488 8576
rect 50356 8430 50384 8570
rect 50252 8424 50304 8430
rect 50252 8366 50304 8372
rect 50344 8424 50396 8430
rect 50344 8366 50396 8372
rect 49792 7880 49844 7886
rect 49792 7822 49844 7828
rect 49332 6792 49384 6798
rect 49330 6760 49332 6769
rect 49516 6792 49568 6798
rect 49384 6760 49386 6769
rect 49516 6734 49568 6740
rect 49330 6695 49386 6704
rect 49332 6384 49384 6390
rect 49792 6384 49844 6390
rect 49332 6326 49384 6332
rect 49620 6332 49792 6338
rect 49620 6326 49844 6332
rect 49344 6089 49372 6326
rect 49620 6310 49832 6326
rect 49516 6248 49568 6254
rect 49514 6216 49516 6225
rect 49568 6216 49570 6225
rect 49620 6186 49648 6310
rect 49514 6151 49570 6160
rect 49608 6180 49660 6186
rect 49608 6122 49660 6128
rect 49792 6180 49844 6186
rect 49792 6122 49844 6128
rect 49330 6080 49386 6089
rect 49330 6015 49386 6024
rect 49422 5944 49478 5953
rect 49422 5879 49424 5888
rect 49476 5879 49478 5888
rect 49424 5850 49476 5856
rect 49238 5808 49294 5817
rect 49238 5743 49294 5752
rect 49252 5710 49280 5743
rect 49804 5710 49832 6122
rect 50264 5914 50292 8366
rect 50448 7954 50476 8570
rect 50436 7948 50488 7954
rect 50436 7890 50488 7896
rect 50448 7274 50476 7890
rect 50436 7268 50488 7274
rect 50436 7210 50488 7216
rect 50540 6440 50568 11494
rect 50632 11286 50660 11562
rect 51092 11558 51120 12718
rect 52564 12374 52592 13806
rect 53024 13462 53052 14418
rect 54024 13864 54076 13870
rect 54024 13806 54076 13812
rect 54576 13864 54628 13870
rect 54576 13806 54628 13812
rect 53564 13796 53616 13802
rect 53564 13738 53616 13744
rect 53932 13796 53984 13802
rect 53932 13738 53984 13744
rect 53012 13456 53064 13462
rect 53012 13398 53064 13404
rect 53104 13388 53156 13394
rect 53104 13330 53156 13336
rect 53380 13388 53432 13394
rect 53380 13330 53432 13336
rect 52736 12708 52788 12714
rect 52736 12650 52788 12656
rect 52552 12368 52604 12374
rect 52552 12310 52604 12316
rect 51862 11996 52158 12016
rect 51918 11994 51942 11996
rect 51998 11994 52022 11996
rect 52078 11994 52102 11996
rect 51940 11942 51942 11994
rect 52004 11942 52016 11994
rect 52078 11942 52080 11994
rect 51918 11940 51942 11942
rect 51998 11940 52022 11942
rect 52078 11940 52102 11942
rect 51862 11920 52158 11940
rect 52000 11824 52052 11830
rect 52000 11766 52052 11772
rect 51632 11688 51684 11694
rect 51632 11630 51684 11636
rect 51080 11552 51132 11558
rect 51080 11494 51132 11500
rect 51540 11348 51592 11354
rect 51540 11290 51592 11296
rect 50620 11280 50672 11286
rect 50620 11222 50672 11228
rect 51552 11150 51580 11290
rect 51540 11144 51592 11150
rect 51540 11086 51592 11092
rect 51356 10532 51408 10538
rect 51356 10474 51408 10480
rect 51368 10130 51396 10474
rect 51448 10464 51500 10470
rect 51448 10406 51500 10412
rect 51356 10124 51408 10130
rect 51356 10066 51408 10072
rect 51264 9512 51316 9518
rect 51264 9454 51316 9460
rect 50804 8288 50856 8294
rect 50804 8230 50856 8236
rect 50816 7886 50844 8230
rect 50804 7880 50856 7886
rect 50804 7822 50856 7828
rect 51276 7818 51304 9454
rect 51460 9042 51488 10406
rect 51552 10062 51580 11086
rect 51540 10056 51592 10062
rect 51540 9998 51592 10004
rect 51552 9518 51580 9998
rect 51540 9512 51592 9518
rect 51540 9454 51592 9460
rect 51448 9036 51500 9042
rect 51448 8978 51500 8984
rect 51356 8968 51408 8974
rect 51356 8910 51408 8916
rect 51368 8566 51396 8910
rect 51356 8560 51408 8566
rect 51356 8502 51408 8508
rect 51460 7954 51488 8978
rect 51448 7948 51500 7954
rect 51448 7890 51500 7896
rect 51264 7812 51316 7818
rect 51264 7754 51316 7760
rect 51552 7342 51580 9454
rect 51540 7336 51592 7342
rect 51540 7278 51592 7284
rect 51356 6928 51408 6934
rect 51262 6896 51318 6905
rect 51356 6870 51408 6876
rect 51262 6831 51264 6840
rect 51316 6831 51318 6840
rect 51264 6802 51316 6808
rect 51264 6656 51316 6662
rect 51264 6598 51316 6604
rect 51276 6497 51304 6598
rect 50448 6412 50568 6440
rect 51262 6488 51318 6497
rect 51262 6423 51318 6432
rect 50252 5908 50304 5914
rect 50252 5850 50304 5856
rect 49884 5840 49936 5846
rect 49884 5782 49936 5788
rect 49240 5704 49292 5710
rect 49240 5646 49292 5652
rect 49792 5704 49844 5710
rect 49792 5646 49844 5652
rect 49804 5166 49832 5646
rect 49896 5522 49924 5782
rect 50448 5778 50476 6412
rect 50710 6352 50766 6361
rect 50528 6316 50580 6322
rect 50710 6287 50766 6296
rect 51170 6352 51226 6361
rect 51170 6287 51172 6296
rect 50528 6258 50580 6264
rect 50540 5914 50568 6258
rect 50620 6248 50672 6254
rect 50620 6190 50672 6196
rect 50528 5908 50580 5914
rect 50528 5850 50580 5856
rect 50632 5846 50660 6190
rect 50724 6118 50752 6287
rect 51224 6287 51226 6296
rect 51172 6258 51224 6264
rect 50712 6112 50764 6118
rect 50712 6054 50764 6060
rect 50620 5840 50672 5846
rect 50620 5782 50672 5788
rect 50436 5772 50488 5778
rect 50436 5714 50488 5720
rect 51264 5772 51316 5778
rect 51264 5714 51316 5720
rect 49896 5494 50016 5522
rect 49608 5160 49660 5166
rect 49608 5102 49660 5108
rect 49792 5160 49844 5166
rect 49792 5102 49844 5108
rect 49056 4684 49108 4690
rect 49056 4626 49108 4632
rect 48780 4616 48832 4622
rect 48780 4558 48832 4564
rect 49424 4616 49476 4622
rect 49424 4558 49476 4564
rect 49436 4214 49464 4558
rect 49424 4208 49476 4214
rect 49424 4150 49476 4156
rect 49516 4072 49568 4078
rect 49620 4026 49648 5102
rect 49988 5030 50016 5494
rect 50068 5296 50120 5302
rect 50068 5238 50120 5244
rect 49976 5024 50028 5030
rect 49976 4966 50028 4972
rect 49700 4276 49752 4282
rect 49700 4218 49752 4224
rect 49568 4020 49648 4026
rect 49516 4014 49648 4020
rect 49528 3998 49648 4014
rect 49620 3618 49648 3998
rect 49712 3738 49740 4218
rect 49884 4072 49936 4078
rect 49884 4014 49936 4020
rect 49896 3738 49924 4014
rect 49700 3732 49752 3738
rect 49700 3674 49752 3680
rect 49884 3732 49936 3738
rect 49884 3674 49936 3680
rect 49620 3602 49740 3618
rect 49620 3596 49752 3602
rect 49620 3590 49700 3596
rect 49700 3538 49752 3544
rect 49988 3398 50016 4966
rect 50080 4078 50108 5238
rect 50804 5228 50856 5234
rect 50804 5170 50856 5176
rect 50540 5098 50752 5114
rect 50436 5092 50488 5098
rect 50436 5034 50488 5040
rect 50540 5092 50764 5098
rect 50540 5086 50712 5092
rect 50448 4826 50476 5034
rect 50540 5030 50568 5086
rect 50712 5034 50764 5040
rect 50528 5024 50580 5030
rect 50528 4966 50580 4972
rect 50436 4820 50488 4826
rect 50436 4762 50488 4768
rect 50816 4758 50844 5170
rect 50804 4752 50856 4758
rect 50804 4694 50856 4700
rect 50436 4616 50488 4622
rect 50436 4558 50488 4564
rect 50068 4072 50120 4078
rect 50068 4014 50120 4020
rect 50448 3534 50476 4558
rect 51276 3534 51304 5714
rect 51368 4282 51396 6870
rect 51644 6390 51672 11630
rect 52012 11218 52040 11766
rect 52368 11552 52420 11558
rect 52368 11494 52420 11500
rect 52000 11212 52052 11218
rect 52000 11154 52052 11160
rect 51862 10908 52158 10928
rect 51918 10906 51942 10908
rect 51998 10906 52022 10908
rect 52078 10906 52102 10908
rect 51940 10854 51942 10906
rect 52004 10854 52016 10906
rect 52078 10854 52080 10906
rect 51918 10852 51942 10854
rect 51998 10852 52022 10854
rect 52078 10852 52102 10854
rect 51862 10832 52158 10852
rect 52380 10674 52408 11494
rect 52368 10668 52420 10674
rect 52368 10610 52420 10616
rect 51724 10056 51776 10062
rect 51724 9998 51776 10004
rect 51736 9450 51764 9998
rect 51862 9820 52158 9840
rect 51918 9818 51942 9820
rect 51998 9818 52022 9820
rect 52078 9818 52102 9820
rect 51940 9766 51942 9818
rect 52004 9766 52016 9818
rect 52078 9766 52080 9818
rect 51918 9764 51942 9766
rect 51998 9764 52022 9766
rect 52078 9764 52102 9766
rect 51862 9744 52158 9764
rect 52748 9636 52776 12650
rect 52920 11892 52972 11898
rect 52920 11834 52972 11840
rect 52932 11665 52960 11834
rect 52918 11656 52974 11665
rect 52918 11591 52974 11600
rect 52932 10606 52960 11591
rect 53116 10810 53144 13330
rect 53196 13320 53248 13326
rect 53196 13262 53248 13268
rect 53208 12850 53236 13262
rect 53196 12844 53248 12850
rect 53196 12786 53248 12792
rect 53208 12442 53236 12786
rect 53196 12436 53248 12442
rect 53196 12378 53248 12384
rect 53196 11688 53248 11694
rect 53196 11630 53248 11636
rect 53208 11354 53236 11630
rect 53196 11348 53248 11354
rect 53196 11290 53248 11296
rect 53104 10804 53156 10810
rect 53104 10746 53156 10752
rect 52920 10600 52972 10606
rect 52920 10542 52972 10548
rect 53196 10532 53248 10538
rect 53196 10474 53248 10480
rect 53208 9926 53236 10474
rect 53196 9920 53248 9926
rect 53196 9862 53248 9868
rect 52656 9608 52776 9636
rect 51724 9444 51776 9450
rect 51724 9386 51776 9392
rect 51724 9036 51776 9042
rect 51724 8978 51776 8984
rect 51736 8022 51764 8978
rect 52184 8900 52236 8906
rect 52184 8842 52236 8848
rect 51862 8732 52158 8752
rect 51918 8730 51942 8732
rect 51998 8730 52022 8732
rect 52078 8730 52102 8732
rect 51940 8678 51942 8730
rect 52004 8678 52016 8730
rect 52078 8678 52080 8730
rect 51918 8676 51942 8678
rect 51998 8676 52022 8678
rect 52078 8676 52102 8678
rect 51862 8656 52158 8676
rect 52196 8430 52224 8842
rect 52184 8424 52236 8430
rect 52184 8366 52236 8372
rect 51724 8016 51776 8022
rect 51724 7958 51776 7964
rect 52460 7948 52512 7954
rect 52460 7890 52512 7896
rect 51862 7644 52158 7664
rect 51918 7642 51942 7644
rect 51998 7642 52022 7644
rect 52078 7642 52102 7644
rect 51940 7590 51942 7642
rect 52004 7590 52016 7642
rect 52078 7590 52080 7642
rect 51918 7588 51942 7590
rect 51998 7588 52022 7590
rect 52078 7588 52102 7590
rect 51862 7568 52158 7588
rect 51724 7336 51776 7342
rect 51724 7278 51776 7284
rect 51632 6384 51684 6390
rect 51632 6326 51684 6332
rect 51448 6248 51500 6254
rect 51448 6190 51500 6196
rect 51460 5370 51488 6190
rect 51540 5840 51592 5846
rect 51540 5782 51592 5788
rect 51552 5370 51580 5782
rect 51448 5364 51500 5370
rect 51448 5306 51500 5312
rect 51540 5364 51592 5370
rect 51540 5306 51592 5312
rect 51736 4690 51764 7278
rect 52368 6792 52420 6798
rect 52472 6769 52500 7890
rect 52552 7336 52604 7342
rect 52552 7278 52604 7284
rect 52564 6934 52592 7278
rect 52552 6928 52604 6934
rect 52552 6870 52604 6876
rect 52368 6734 52420 6740
rect 52458 6760 52514 6769
rect 52184 6724 52236 6730
rect 52184 6666 52236 6672
rect 51862 6556 52158 6576
rect 51918 6554 51942 6556
rect 51998 6554 52022 6556
rect 52078 6554 52102 6556
rect 51940 6502 51942 6554
rect 52004 6502 52016 6554
rect 52078 6502 52080 6554
rect 51918 6500 51942 6502
rect 51998 6500 52022 6502
rect 52078 6500 52102 6502
rect 51862 6480 52158 6500
rect 52196 6390 52224 6666
rect 52184 6384 52236 6390
rect 52184 6326 52236 6332
rect 52274 6216 52330 6225
rect 52274 6151 52330 6160
rect 52184 6112 52236 6118
rect 52184 6054 52236 6060
rect 52196 5817 52224 6054
rect 52182 5808 52238 5817
rect 52092 5772 52144 5778
rect 52182 5743 52238 5752
rect 52092 5714 52144 5720
rect 52104 5642 52132 5714
rect 52092 5636 52144 5642
rect 52092 5578 52144 5584
rect 52288 5574 52316 6151
rect 52380 5642 52408 6734
rect 52458 6695 52514 6704
rect 52656 6236 52684 9608
rect 52736 9512 52788 9518
rect 52736 9454 52788 9460
rect 52748 8634 52776 9454
rect 52920 9376 52972 9382
rect 52920 9318 52972 9324
rect 52932 9110 52960 9318
rect 52920 9104 52972 9110
rect 52920 9046 52972 9052
rect 53208 8974 53236 9862
rect 53196 8968 53248 8974
rect 53196 8910 53248 8916
rect 52736 8628 52788 8634
rect 52736 8570 52788 8576
rect 53196 8424 53248 8430
rect 53196 8366 53248 8372
rect 53104 7880 53156 7886
rect 53104 7822 53156 7828
rect 52920 6656 52972 6662
rect 52918 6624 52920 6633
rect 53012 6656 53064 6662
rect 52972 6624 52974 6633
rect 53012 6598 53064 6604
rect 52918 6559 52974 6568
rect 53024 6458 53052 6598
rect 53012 6452 53064 6458
rect 53012 6394 53064 6400
rect 52828 6248 52880 6254
rect 52656 6208 52828 6236
rect 52828 6190 52880 6196
rect 52840 5914 52868 6190
rect 53012 6180 53064 6186
rect 53012 6122 53064 6128
rect 52460 5908 52512 5914
rect 52460 5850 52512 5856
rect 52828 5908 52880 5914
rect 52828 5850 52880 5856
rect 52368 5636 52420 5642
rect 52368 5578 52420 5584
rect 52276 5568 52328 5574
rect 52276 5510 52328 5516
rect 51862 5468 52158 5488
rect 51918 5466 51942 5468
rect 51998 5466 52022 5468
rect 52078 5466 52102 5468
rect 51940 5414 51942 5466
rect 52004 5414 52016 5466
rect 52078 5414 52080 5466
rect 51918 5412 51942 5414
rect 51998 5412 52022 5414
rect 52078 5412 52102 5414
rect 51862 5392 52158 5412
rect 52472 4690 52500 5850
rect 53024 5370 53052 6122
rect 53012 5364 53064 5370
rect 53012 5306 53064 5312
rect 51724 4684 51776 4690
rect 51724 4626 51776 4632
rect 52460 4684 52512 4690
rect 52460 4626 52512 4632
rect 51356 4276 51408 4282
rect 51356 4218 51408 4224
rect 51736 4146 51764 4626
rect 52276 4616 52328 4622
rect 52276 4558 52328 4564
rect 51862 4380 52158 4400
rect 51918 4378 51942 4380
rect 51998 4378 52022 4380
rect 52078 4378 52102 4380
rect 51940 4326 51942 4378
rect 52004 4326 52016 4378
rect 52078 4326 52080 4378
rect 51918 4324 51942 4326
rect 51998 4324 52022 4326
rect 52078 4324 52102 4326
rect 51862 4304 52158 4324
rect 52288 4282 52316 4558
rect 52276 4276 52328 4282
rect 52276 4218 52328 4224
rect 51724 4140 51776 4146
rect 51724 4082 51776 4088
rect 51632 3936 51684 3942
rect 51632 3878 51684 3884
rect 51644 3602 51672 3878
rect 53116 3641 53144 7822
rect 53208 7206 53236 8366
rect 53196 7200 53248 7206
rect 53196 7142 53248 7148
rect 53208 6934 53236 7142
rect 53196 6928 53248 6934
rect 53196 6870 53248 6876
rect 53288 6792 53340 6798
rect 53288 6734 53340 6740
rect 53300 6254 53328 6734
rect 53288 6248 53340 6254
rect 53288 6190 53340 6196
rect 53392 5778 53420 13330
rect 53576 13326 53604 13738
rect 53944 13530 53972 13738
rect 53932 13524 53984 13530
rect 53932 13466 53984 13472
rect 53564 13320 53616 13326
rect 53564 13262 53616 13268
rect 53576 12850 53604 13262
rect 54036 12986 54064 13806
rect 54024 12980 54076 12986
rect 54024 12922 54076 12928
rect 53564 12844 53616 12850
rect 53564 12786 53616 12792
rect 53576 12306 53604 12786
rect 54588 12374 54616 13806
rect 54680 13462 54708 15370
rect 55324 15026 55352 16594
rect 55496 15360 55548 15366
rect 55496 15302 55548 15308
rect 55312 15020 55364 15026
rect 55312 14962 55364 14968
rect 55036 14952 55088 14958
rect 55036 14894 55088 14900
rect 55220 14952 55272 14958
rect 55220 14894 55272 14900
rect 54852 14408 54904 14414
rect 54852 14350 54904 14356
rect 54864 13938 54892 14350
rect 55048 14074 55076 14894
rect 55036 14068 55088 14074
rect 55036 14010 55088 14016
rect 54852 13932 54904 13938
rect 54852 13874 54904 13880
rect 54668 13456 54720 13462
rect 54668 13398 54720 13404
rect 55232 12986 55260 14894
rect 55324 14482 55352 14962
rect 55312 14476 55364 14482
rect 55312 14418 55364 14424
rect 55508 13870 55536 15302
rect 55600 15162 55628 16594
rect 55864 15904 55916 15910
rect 55864 15846 55916 15852
rect 55588 15156 55640 15162
rect 55588 15098 55640 15104
rect 55876 14890 55904 15846
rect 55864 14884 55916 14890
rect 55864 14826 55916 14832
rect 56520 14550 56548 18835
rect 58452 16590 58480 18835
rect 57060 16584 57112 16590
rect 57060 16526 57112 16532
rect 58440 16584 58492 16590
rect 58440 16526 58492 16532
rect 57072 16046 57100 16526
rect 57060 16040 57112 16046
rect 57060 15982 57112 15988
rect 60384 15638 60412 18835
rect 62316 16114 62344 18835
rect 62304 16108 62356 16114
rect 62304 16050 62356 16056
rect 58716 15632 58768 15638
rect 58716 15574 58768 15580
rect 60372 15632 60424 15638
rect 60372 15574 60424 15580
rect 58728 14550 58756 15574
rect 56508 14544 56560 14550
rect 56508 14486 56560 14492
rect 58716 14544 58768 14550
rect 58716 14486 58768 14492
rect 56416 14408 56468 14414
rect 56416 14350 56468 14356
rect 55496 13864 55548 13870
rect 55496 13806 55548 13812
rect 55220 12980 55272 12986
rect 55220 12922 55272 12928
rect 56428 12850 56456 14350
rect 56520 13394 56548 14486
rect 57336 14408 57388 14414
rect 57336 14350 57388 14356
rect 57348 13938 57376 14350
rect 57336 13932 57388 13938
rect 57336 13874 57388 13880
rect 56508 13388 56560 13394
rect 56508 13330 56560 13336
rect 55036 12844 55088 12850
rect 55036 12786 55088 12792
rect 56416 12844 56468 12850
rect 56416 12786 56468 12792
rect 55048 12442 55076 12786
rect 55312 12776 55364 12782
rect 55312 12718 55364 12724
rect 55772 12776 55824 12782
rect 55772 12718 55824 12724
rect 58440 12776 58492 12782
rect 58440 12718 58492 12724
rect 55036 12436 55088 12442
rect 55036 12378 55088 12384
rect 54576 12368 54628 12374
rect 54576 12310 54628 12316
rect 55048 12306 55076 12378
rect 53472 12300 53524 12306
rect 53472 12242 53524 12248
rect 53564 12300 53616 12306
rect 53564 12242 53616 12248
rect 55036 12300 55088 12306
rect 55036 12242 55088 12248
rect 53484 5846 53512 12242
rect 53748 12232 53800 12238
rect 53748 12174 53800 12180
rect 53760 11286 53788 12174
rect 55220 12164 55272 12170
rect 55220 12106 55272 12112
rect 55232 12050 55260 12106
rect 55140 12022 55260 12050
rect 54668 11552 54720 11558
rect 54668 11494 54720 11500
rect 53748 11280 53800 11286
rect 53748 11222 53800 11228
rect 54680 11218 54708 11494
rect 54668 11212 54720 11218
rect 54668 11154 54720 11160
rect 54576 11144 54628 11150
rect 54576 11086 54628 11092
rect 54588 11014 54616 11086
rect 54576 11008 54628 11014
rect 54576 10950 54628 10956
rect 54300 10600 54352 10606
rect 54300 10542 54352 10548
rect 54312 9382 54340 10542
rect 54588 10062 54616 10950
rect 54760 10464 54812 10470
rect 54760 10406 54812 10412
rect 54668 10124 54720 10130
rect 54668 10066 54720 10072
rect 54576 10056 54628 10062
rect 54576 9998 54628 10004
rect 54680 9586 54708 10066
rect 54668 9580 54720 9586
rect 54668 9522 54720 9528
rect 54300 9376 54352 9382
rect 54300 9318 54352 9324
rect 54680 9110 54708 9522
rect 54772 9450 54800 10406
rect 54852 9920 54904 9926
rect 54852 9862 54904 9868
rect 54864 9654 54892 9862
rect 54852 9648 54904 9654
rect 54852 9590 54904 9596
rect 54864 9518 54892 9590
rect 54852 9512 54904 9518
rect 54852 9454 54904 9460
rect 54760 9444 54812 9450
rect 54760 9386 54812 9392
rect 54668 9104 54720 9110
rect 54668 9046 54720 9052
rect 54772 9042 54800 9386
rect 53656 9036 53708 9042
rect 53656 8978 53708 8984
rect 54760 9036 54812 9042
rect 54760 8978 54812 8984
rect 53668 8430 53696 8978
rect 54864 8974 54892 9454
rect 54944 9036 54996 9042
rect 54944 8978 54996 8984
rect 54852 8968 54904 8974
rect 54852 8910 54904 8916
rect 54956 8498 54984 8978
rect 55036 8900 55088 8906
rect 55036 8842 55088 8848
rect 55048 8634 55076 8842
rect 55036 8628 55088 8634
rect 55036 8570 55088 8576
rect 54944 8492 54996 8498
rect 54944 8434 54996 8440
rect 53656 8424 53708 8430
rect 53654 8392 53656 8401
rect 53708 8392 53710 8401
rect 53654 8327 53710 8336
rect 55048 7954 55076 8570
rect 55036 7948 55088 7954
rect 55036 7890 55088 7896
rect 53748 7812 53800 7818
rect 53748 7754 53800 7760
rect 54852 7812 54904 7818
rect 54852 7754 54904 7760
rect 53656 6928 53708 6934
rect 53656 6870 53708 6876
rect 53668 6474 53696 6870
rect 53760 6798 53788 7754
rect 54760 7404 54812 7410
rect 54760 7346 54812 7352
rect 54772 7274 54800 7346
rect 53932 7268 53984 7274
rect 53932 7210 53984 7216
rect 54760 7268 54812 7274
rect 54760 7210 54812 7216
rect 53840 6860 53892 6866
rect 53840 6802 53892 6808
rect 53748 6792 53800 6798
rect 53748 6734 53800 6740
rect 53746 6624 53802 6633
rect 53746 6559 53802 6568
rect 53576 6458 53696 6474
rect 53760 6458 53788 6559
rect 53564 6452 53696 6458
rect 53616 6446 53696 6452
rect 53748 6452 53800 6458
rect 53564 6394 53616 6400
rect 53748 6394 53800 6400
rect 53746 6352 53802 6361
rect 53564 6316 53616 6322
rect 53746 6287 53802 6296
rect 53564 6258 53616 6264
rect 53576 5953 53604 6258
rect 53760 6186 53788 6287
rect 53748 6180 53800 6186
rect 53748 6122 53800 6128
rect 53562 5944 53618 5953
rect 53562 5879 53618 5888
rect 53472 5840 53524 5846
rect 53472 5782 53524 5788
rect 53380 5772 53432 5778
rect 53380 5714 53432 5720
rect 53392 5234 53420 5714
rect 53484 5302 53512 5782
rect 53852 5642 53880 6802
rect 53944 6361 53972 7210
rect 54022 6896 54078 6905
rect 54772 6866 54800 7210
rect 54022 6831 54078 6840
rect 54760 6860 54812 6866
rect 54036 6662 54064 6831
rect 54760 6802 54812 6808
rect 54024 6656 54076 6662
rect 54024 6598 54076 6604
rect 53930 6352 53986 6361
rect 53930 6287 53932 6296
rect 53984 6287 53986 6296
rect 54668 6316 54720 6322
rect 53932 6258 53984 6264
rect 54668 6258 54720 6264
rect 53944 6227 53972 6258
rect 54484 6248 54536 6254
rect 54576 6248 54628 6254
rect 54536 6208 54576 6236
rect 54484 6190 54536 6196
rect 54576 6190 54628 6196
rect 54680 6089 54708 6258
rect 54666 6080 54722 6089
rect 54666 6015 54722 6024
rect 54772 5710 54800 6802
rect 54760 5704 54812 5710
rect 54760 5646 54812 5652
rect 53840 5636 53892 5642
rect 53840 5578 53892 5584
rect 54392 5636 54444 5642
rect 54392 5578 54444 5584
rect 53472 5296 53524 5302
rect 53472 5238 53524 5244
rect 53380 5228 53432 5234
rect 53380 5170 53432 5176
rect 53748 5160 53800 5166
rect 53748 5102 53800 5108
rect 53472 4072 53524 4078
rect 53472 4014 53524 4020
rect 53102 3632 53158 3641
rect 51632 3596 51684 3602
rect 53102 3567 53158 3576
rect 51632 3538 51684 3544
rect 50436 3528 50488 3534
rect 50436 3470 50488 3476
rect 51264 3528 51316 3534
rect 51264 3470 51316 3476
rect 52184 3528 52236 3534
rect 52184 3470 52236 3476
rect 53196 3528 53248 3534
rect 53196 3470 53248 3476
rect 50620 3460 50672 3466
rect 50620 3402 50672 3408
rect 49976 3392 50028 3398
rect 49976 3334 50028 3340
rect 48686 3224 48742 3233
rect 48686 3159 48742 3168
rect 49988 2990 50016 3334
rect 49792 2984 49844 2990
rect 49792 2926 49844 2932
rect 49976 2984 50028 2990
rect 49976 2926 50028 2932
rect 49804 2854 49832 2926
rect 49792 2848 49844 2854
rect 49792 2790 49844 2796
rect 48596 2644 48648 2650
rect 48596 2586 48648 2592
rect 41052 2508 41104 2514
rect 41052 2450 41104 2456
rect 41328 2508 41380 2514
rect 41328 2450 41380 2456
rect 44548 2508 44600 2514
rect 44548 2450 44600 2456
rect 48044 2508 48096 2514
rect 48044 2450 48096 2456
rect 48504 2508 48556 2514
rect 48504 2450 48556 2456
rect 40500 2100 40552 2106
rect 40500 2042 40552 2048
rect 41064 800 41092 2450
rect 43720 2440 43772 2446
rect 43720 2382 43772 2388
rect 41972 2372 42024 2378
rect 41972 2314 42024 2320
rect 41984 800 42012 2314
rect 42800 2304 42852 2310
rect 42800 2246 42852 2252
rect 42892 2304 42944 2310
rect 42892 2246 42944 2252
rect 42812 2038 42840 2246
rect 42800 2032 42852 2038
rect 42800 1974 42852 1980
rect 42904 1170 42932 2246
rect 42812 1142 42932 1170
rect 42812 800 42840 1142
rect 43732 800 43760 2382
rect 44560 800 44588 2450
rect 47124 2440 47176 2446
rect 47124 2382 47176 2388
rect 45468 2372 45520 2378
rect 45468 2314 45520 2320
rect 46296 2372 46348 2378
rect 46296 2314 46348 2320
rect 45480 800 45508 2314
rect 46308 800 46336 2314
rect 47136 800 47164 2382
rect 48056 800 48084 2450
rect 49792 2440 49844 2446
rect 49792 2382 49844 2388
rect 48872 2304 48924 2310
rect 48872 2246 48924 2252
rect 48884 800 48912 2246
rect 49804 800 49832 2382
rect 50632 800 50660 3402
rect 51276 3194 51304 3470
rect 51540 3392 51592 3398
rect 51540 3334 51592 3340
rect 51264 3188 51316 3194
rect 51264 3130 51316 3136
rect 51552 800 51580 3334
rect 51862 3292 52158 3312
rect 51918 3290 51942 3292
rect 51998 3290 52022 3292
rect 52078 3290 52102 3292
rect 51940 3238 51942 3290
rect 52004 3238 52016 3290
rect 52078 3238 52080 3290
rect 51918 3236 51942 3238
rect 51998 3236 52022 3238
rect 52078 3236 52102 3238
rect 51862 3216 52158 3236
rect 52196 3058 52224 3470
rect 52460 3188 52512 3194
rect 52460 3130 52512 3136
rect 52184 3052 52236 3058
rect 52184 2994 52236 3000
rect 52472 2961 52500 3130
rect 52458 2952 52514 2961
rect 52458 2887 52514 2896
rect 52368 2304 52420 2310
rect 52368 2246 52420 2252
rect 51862 2204 52158 2224
rect 51918 2202 51942 2204
rect 51998 2202 52022 2204
rect 52078 2202 52102 2204
rect 51940 2150 51942 2202
rect 52004 2150 52016 2202
rect 52078 2150 52080 2202
rect 51918 2148 51942 2150
rect 51998 2148 52022 2150
rect 52078 2148 52102 2150
rect 51862 2128 52158 2148
rect 52380 800 52408 2246
rect 53208 800 53236 3470
rect 53484 3194 53512 4014
rect 53760 3942 53788 5102
rect 54024 4140 54076 4146
rect 54024 4082 54076 4088
rect 53748 3936 53800 3942
rect 53748 3878 53800 3884
rect 53564 3392 53616 3398
rect 53564 3334 53616 3340
rect 53576 3194 53604 3334
rect 53472 3188 53524 3194
rect 53472 3130 53524 3136
rect 53564 3188 53616 3194
rect 53564 3130 53616 3136
rect 53760 2990 53788 3878
rect 54036 3641 54064 4082
rect 54022 3632 54078 3641
rect 54022 3567 54078 3576
rect 54036 2990 54064 3567
rect 54404 2990 54432 5578
rect 54864 5166 54892 7754
rect 55140 6361 55168 12022
rect 55324 11762 55352 12718
rect 55784 12306 55812 12718
rect 56140 12708 56192 12714
rect 56140 12650 56192 12656
rect 55864 12368 55916 12374
rect 55864 12310 55916 12316
rect 55772 12300 55824 12306
rect 55772 12242 55824 12248
rect 55876 11898 55904 12310
rect 56048 12232 56100 12238
rect 56048 12174 56100 12180
rect 55864 11892 55916 11898
rect 55864 11834 55916 11840
rect 56060 11830 56088 12174
rect 56048 11824 56100 11830
rect 56048 11766 56100 11772
rect 55312 11756 55364 11762
rect 55312 11698 55364 11704
rect 56060 10606 56088 11766
rect 55404 10600 55456 10606
rect 55404 10542 55456 10548
rect 56048 10600 56100 10606
rect 56048 10542 56100 10548
rect 55312 8832 55364 8838
rect 55312 8774 55364 8780
rect 55220 8560 55272 8566
rect 55220 8502 55272 8508
rect 55232 8090 55260 8502
rect 55220 8084 55272 8090
rect 55220 8026 55272 8032
rect 55324 7954 55352 8774
rect 55312 7948 55364 7954
rect 55312 7890 55364 7896
rect 55416 7886 55444 10542
rect 55772 10532 55824 10538
rect 55772 10474 55824 10480
rect 55784 10198 55812 10474
rect 55772 10192 55824 10198
rect 55772 10134 55824 10140
rect 55772 9444 55824 9450
rect 55772 9386 55824 9392
rect 55784 8022 55812 9386
rect 55862 8528 55918 8537
rect 55862 8463 55918 8472
rect 55876 8430 55904 8463
rect 55864 8424 55916 8430
rect 55864 8366 55916 8372
rect 55772 8016 55824 8022
rect 55772 7958 55824 7964
rect 55404 7880 55456 7886
rect 55404 7822 55456 7828
rect 55680 7880 55732 7886
rect 55680 7822 55732 7828
rect 55126 6352 55182 6361
rect 55126 6287 55182 6296
rect 55140 6254 55168 6287
rect 55128 6248 55180 6254
rect 55128 6190 55180 6196
rect 55404 6248 55456 6254
rect 55404 6190 55456 6196
rect 55416 5846 55444 6190
rect 55404 5840 55456 5846
rect 55404 5782 55456 5788
rect 55312 5364 55364 5370
rect 55312 5306 55364 5312
rect 54852 5160 54904 5166
rect 54852 5102 54904 5108
rect 55324 4434 55352 5306
rect 55404 5092 55456 5098
rect 55404 5034 55456 5040
rect 55416 4554 55444 5034
rect 55404 4548 55456 4554
rect 55404 4490 55456 4496
rect 55692 4486 55720 7822
rect 55784 7342 55812 7958
rect 55772 7336 55824 7342
rect 55772 7278 55824 7284
rect 55864 7336 55916 7342
rect 55864 7278 55916 7284
rect 55680 4480 55732 4486
rect 55324 4406 55444 4434
rect 55680 4422 55732 4428
rect 55312 4140 55364 4146
rect 55312 4082 55364 4088
rect 55324 3602 55352 4082
rect 55416 4078 55444 4406
rect 55404 4072 55456 4078
rect 55404 4014 55456 4020
rect 55312 3596 55364 3602
rect 55312 3538 55364 3544
rect 54576 3528 54628 3534
rect 54576 3470 54628 3476
rect 54588 2990 54616 3470
rect 55416 3058 55444 4014
rect 55588 3936 55640 3942
rect 55588 3878 55640 3884
rect 55600 3534 55628 3878
rect 55692 3602 55720 4422
rect 55876 4078 55904 7278
rect 56152 6866 56180 12650
rect 58164 12300 58216 12306
rect 58164 12242 58216 12248
rect 56232 12096 56284 12102
rect 56232 12038 56284 12044
rect 56244 11694 56272 12038
rect 56784 11756 56836 11762
rect 56784 11698 56836 11704
rect 56232 11688 56284 11694
rect 56600 11688 56652 11694
rect 56284 11636 56364 11642
rect 56232 11630 56364 11636
rect 56600 11630 56652 11636
rect 56244 11614 56364 11630
rect 56232 11552 56284 11558
rect 56232 11494 56284 11500
rect 56244 11082 56272 11494
rect 56336 11354 56364 11614
rect 56324 11348 56376 11354
rect 56324 11290 56376 11296
rect 56612 11150 56640 11630
rect 56692 11620 56744 11626
rect 56692 11562 56744 11568
rect 56704 11218 56732 11562
rect 56692 11212 56744 11218
rect 56692 11154 56744 11160
rect 56600 11144 56652 11150
rect 56600 11086 56652 11092
rect 56232 11076 56284 11082
rect 56232 11018 56284 11024
rect 56244 10606 56272 11018
rect 56232 10600 56284 10606
rect 56232 10542 56284 10548
rect 56612 9994 56640 11086
rect 56796 10742 56824 11698
rect 57336 11688 57388 11694
rect 57336 11630 57388 11636
rect 57348 11014 57376 11630
rect 57336 11008 57388 11014
rect 57336 10950 57388 10956
rect 56784 10736 56836 10742
rect 56784 10678 56836 10684
rect 57348 10674 57376 10950
rect 57336 10668 57388 10674
rect 57336 10610 57388 10616
rect 57348 10062 57376 10610
rect 57336 10056 57388 10062
rect 57336 9998 57388 10004
rect 58072 10056 58124 10062
rect 58072 9998 58124 10004
rect 56600 9988 56652 9994
rect 56600 9930 56652 9936
rect 57348 9518 57376 9998
rect 57336 9512 57388 9518
rect 57336 9454 57388 9460
rect 57980 9512 58032 9518
rect 57980 9454 58032 9460
rect 57058 9072 57114 9081
rect 56692 9036 56744 9042
rect 57058 9007 57060 9016
rect 56692 8978 56744 8984
rect 57112 9007 57114 9016
rect 57244 9036 57296 9042
rect 57060 8978 57112 8984
rect 57244 8978 57296 8984
rect 56704 8945 56732 8978
rect 56690 8936 56746 8945
rect 56690 8871 56746 8880
rect 56876 8900 56928 8906
rect 56876 8842 56928 8848
rect 56324 8424 56376 8430
rect 56324 8366 56376 8372
rect 56140 6860 56192 6866
rect 56140 6802 56192 6808
rect 56152 5930 56180 6802
rect 56232 6792 56284 6798
rect 56232 6734 56284 6740
rect 56244 6118 56272 6734
rect 56232 6112 56284 6118
rect 56232 6054 56284 6060
rect 56152 5902 56272 5930
rect 56244 5710 56272 5902
rect 56232 5704 56284 5710
rect 56232 5646 56284 5652
rect 56336 5574 56364 8366
rect 56888 8362 56916 8842
rect 56876 8356 56928 8362
rect 56876 8298 56928 8304
rect 56968 8356 57020 8362
rect 56968 8298 57020 8304
rect 56980 7954 57008 8298
rect 57256 8090 57284 8978
rect 57244 8084 57296 8090
rect 57244 8026 57296 8032
rect 57242 7984 57298 7993
rect 56968 7948 57020 7954
rect 57992 7970 58020 9454
rect 58084 9110 58112 9998
rect 58072 9104 58124 9110
rect 58072 9046 58124 9052
rect 57992 7942 58112 7970
rect 57242 7919 57298 7928
rect 56968 7890 57020 7896
rect 56980 7410 57008 7890
rect 57256 7886 57284 7919
rect 57244 7880 57296 7886
rect 57244 7822 57296 7828
rect 57980 7880 58032 7886
rect 57980 7822 58032 7828
rect 56968 7404 57020 7410
rect 56968 7346 57020 7352
rect 56968 7200 57020 7206
rect 56968 7142 57020 7148
rect 56980 6866 57008 7142
rect 57992 6866 58020 7822
rect 58084 7410 58112 7942
rect 58072 7404 58124 7410
rect 58072 7346 58124 7352
rect 56692 6860 56744 6866
rect 56692 6802 56744 6808
rect 56968 6860 57020 6866
rect 56968 6802 57020 6808
rect 57980 6860 58032 6866
rect 57980 6802 58032 6808
rect 56704 6390 56732 6802
rect 58176 6458 58204 12242
rect 58452 12170 58480 12718
rect 59728 12640 59780 12646
rect 59728 12582 59780 12588
rect 59740 12306 59768 12582
rect 59728 12300 59780 12306
rect 59728 12242 59780 12248
rect 59084 12232 59136 12238
rect 59084 12174 59136 12180
rect 58440 12164 58492 12170
rect 58440 12106 58492 12112
rect 59096 11354 59124 12174
rect 60464 11892 60516 11898
rect 60464 11834 60516 11840
rect 59084 11348 59136 11354
rect 59084 11290 59136 11296
rect 58716 10464 58768 10470
rect 58716 10406 58768 10412
rect 58728 10130 58756 10406
rect 59360 10260 59412 10266
rect 59360 10202 59412 10208
rect 58716 10124 58768 10130
rect 58716 10066 58768 10072
rect 58532 9920 58584 9926
rect 58532 9862 58584 9868
rect 58348 9512 58400 9518
rect 58348 9454 58400 9460
rect 58360 9178 58388 9454
rect 58348 9172 58400 9178
rect 58348 9114 58400 9120
rect 58544 8634 58572 9862
rect 58716 9036 58768 9042
rect 58716 8978 58768 8984
rect 59268 9036 59320 9042
rect 59268 8978 59320 8984
rect 58728 8945 58756 8978
rect 58808 8968 58860 8974
rect 58714 8936 58770 8945
rect 58808 8910 58860 8916
rect 59176 8968 59228 8974
rect 59176 8910 59228 8916
rect 58714 8871 58770 8880
rect 58532 8628 58584 8634
rect 58532 8570 58584 8576
rect 58544 8430 58572 8570
rect 58532 8424 58584 8430
rect 58532 8366 58584 8372
rect 58348 7744 58400 7750
rect 58348 7686 58400 7692
rect 58164 6452 58216 6458
rect 58164 6394 58216 6400
rect 56692 6384 56744 6390
rect 56692 6326 56744 6332
rect 58072 6180 58124 6186
rect 58072 6122 58124 6128
rect 57796 6112 57848 6118
rect 57796 6054 57848 6060
rect 56508 5908 56560 5914
rect 56508 5850 56560 5856
rect 57520 5908 57572 5914
rect 57520 5850 57572 5856
rect 56324 5568 56376 5574
rect 56324 5510 56376 5516
rect 56336 4690 56364 5510
rect 56520 5166 56548 5850
rect 57532 5710 57560 5850
rect 57808 5778 57836 6054
rect 57796 5772 57848 5778
rect 57796 5714 57848 5720
rect 57520 5704 57572 5710
rect 57520 5646 57572 5652
rect 57532 5370 57560 5646
rect 57704 5636 57756 5642
rect 57704 5578 57756 5584
rect 57520 5364 57572 5370
rect 57520 5306 57572 5312
rect 56508 5160 56560 5166
rect 56508 5102 56560 5108
rect 57612 4752 57664 4758
rect 57612 4694 57664 4700
rect 56324 4684 56376 4690
rect 56324 4626 56376 4632
rect 56508 4684 56560 4690
rect 56508 4626 56560 4632
rect 55864 4072 55916 4078
rect 55864 4014 55916 4020
rect 55956 4072 56008 4078
rect 56520 4049 56548 4626
rect 56692 4548 56744 4554
rect 56692 4490 56744 4496
rect 56704 4146 56732 4490
rect 56692 4140 56744 4146
rect 56692 4082 56744 4088
rect 55956 4014 56008 4020
rect 56506 4040 56562 4049
rect 55968 3942 55996 4014
rect 56506 3975 56562 3984
rect 55956 3936 56008 3942
rect 55956 3878 56008 3884
rect 57624 3738 57652 4694
rect 57716 3942 57744 5578
rect 57808 4078 57836 5714
rect 58084 5234 58112 6122
rect 58360 5574 58388 7686
rect 58440 7404 58492 7410
rect 58440 7346 58492 7352
rect 58348 5568 58400 5574
rect 58348 5510 58400 5516
rect 57980 5228 58032 5234
rect 57980 5170 58032 5176
rect 58072 5228 58124 5234
rect 58072 5170 58124 5176
rect 57992 4622 58020 5170
rect 58452 5166 58480 7346
rect 58624 7336 58676 7342
rect 58624 7278 58676 7284
rect 58636 6934 58664 7278
rect 58624 6928 58676 6934
rect 58624 6870 58676 6876
rect 58728 6866 58756 8871
rect 58820 8566 58848 8910
rect 58808 8560 58860 8566
rect 58808 8502 58860 8508
rect 59188 8498 59216 8910
rect 59176 8492 59228 8498
rect 59176 8434 59228 8440
rect 59280 8430 59308 8978
rect 59268 8424 59320 8430
rect 59268 8366 59320 8372
rect 59268 8016 59320 8022
rect 59268 7958 59320 7964
rect 58808 7744 58860 7750
rect 58808 7686 58860 7692
rect 58820 6866 58848 7686
rect 58716 6860 58768 6866
rect 58716 6802 58768 6808
rect 58808 6860 58860 6866
rect 58808 6802 58860 6808
rect 59280 6730 59308 7958
rect 59372 6934 59400 10202
rect 60188 9376 60240 9382
rect 60188 9318 60240 9324
rect 60200 9042 60228 9318
rect 60188 9036 60240 9042
rect 60188 8978 60240 8984
rect 60280 7948 60332 7954
rect 60280 7890 60332 7896
rect 59452 7880 59504 7886
rect 59452 7822 59504 7828
rect 59360 6928 59412 6934
rect 59360 6870 59412 6876
rect 59268 6724 59320 6730
rect 59268 6666 59320 6672
rect 59280 6322 59308 6666
rect 59268 6316 59320 6322
rect 59268 6258 59320 6264
rect 58716 6248 58768 6254
rect 58716 6190 58768 6196
rect 58808 6248 58860 6254
rect 58808 6190 58860 6196
rect 59176 6248 59228 6254
rect 59176 6190 59228 6196
rect 58624 5568 58676 5574
rect 58624 5510 58676 5516
rect 58440 5160 58492 5166
rect 58492 5108 58572 5114
rect 58440 5102 58572 5108
rect 58452 5086 58572 5102
rect 57980 4616 58032 4622
rect 57980 4558 58032 4564
rect 57796 4072 57848 4078
rect 57796 4014 57848 4020
rect 57992 3942 58020 4558
rect 58440 4548 58492 4554
rect 58440 4490 58492 4496
rect 57704 3936 57756 3942
rect 57704 3878 57756 3884
rect 57980 3936 58032 3942
rect 57980 3878 58032 3884
rect 57612 3732 57664 3738
rect 57612 3674 57664 3680
rect 55864 3664 55916 3670
rect 55864 3606 55916 3612
rect 56874 3632 56930 3641
rect 55680 3596 55732 3602
rect 55680 3538 55732 3544
rect 55588 3528 55640 3534
rect 55588 3470 55640 3476
rect 55772 3528 55824 3534
rect 55772 3470 55824 3476
rect 55600 3097 55628 3470
rect 55586 3088 55642 3097
rect 55404 3052 55456 3058
rect 55586 3023 55642 3032
rect 55404 2994 55456 3000
rect 53748 2984 53800 2990
rect 53748 2926 53800 2932
rect 54024 2984 54076 2990
rect 54024 2926 54076 2932
rect 54392 2984 54444 2990
rect 54392 2926 54444 2932
rect 54576 2984 54628 2990
rect 54576 2926 54628 2932
rect 54668 2984 54720 2990
rect 55588 2984 55640 2990
rect 54668 2926 54720 2932
rect 55586 2952 55588 2961
rect 55784 2972 55812 3470
rect 55640 2952 55812 2972
rect 55642 2944 55812 2952
rect 54680 2854 54708 2926
rect 55586 2887 55642 2896
rect 54668 2848 54720 2854
rect 54668 2790 54720 2796
rect 54944 2508 54996 2514
rect 54944 2450 54996 2456
rect 54116 2304 54168 2310
rect 54116 2246 54168 2252
rect 54128 800 54156 2246
rect 54956 800 54984 2450
rect 55876 800 55904 3606
rect 56784 3596 56836 3602
rect 56874 3567 56876 3576
rect 56784 3538 56836 3544
rect 56928 3567 56930 3576
rect 56876 3538 56928 3544
rect 56692 2984 56744 2990
rect 56692 2926 56744 2932
rect 56704 800 56732 2926
rect 56796 2922 56824 3538
rect 58452 3534 58480 4490
rect 58544 4078 58572 5086
rect 58636 4826 58664 5510
rect 58624 4820 58676 4826
rect 58624 4762 58676 4768
rect 58532 4072 58584 4078
rect 58532 4014 58584 4020
rect 58728 3602 58756 6190
rect 58820 5574 58848 6190
rect 59188 5846 59216 6190
rect 59176 5840 59228 5846
rect 59176 5782 59228 5788
rect 58808 5568 58860 5574
rect 58808 5510 58860 5516
rect 58808 4820 58860 4826
rect 58808 4762 58860 4768
rect 58820 4690 58848 4762
rect 58808 4684 58860 4690
rect 58808 4626 58860 4632
rect 58820 4162 58848 4626
rect 58820 4134 58940 4162
rect 59464 4146 59492 7822
rect 59912 7200 59964 7206
rect 59912 7142 59964 7148
rect 59924 6866 59952 7142
rect 60292 6866 60320 7890
rect 60476 7750 60504 11834
rect 60464 7744 60516 7750
rect 60464 7686 60516 7692
rect 59912 6860 59964 6866
rect 59912 6802 59964 6808
rect 60280 6860 60332 6866
rect 60280 6802 60332 6808
rect 59544 6792 59596 6798
rect 59544 6734 59596 6740
rect 60188 6792 60240 6798
rect 60188 6734 60240 6740
rect 59556 6322 59584 6734
rect 59544 6316 59596 6322
rect 59544 6258 59596 6264
rect 60200 4758 60228 6734
rect 60292 6662 60320 6802
rect 60280 6656 60332 6662
rect 60280 6598 60332 6604
rect 60188 4752 60240 4758
rect 60188 4694 60240 4700
rect 58808 4072 58860 4078
rect 58808 4014 58860 4020
rect 58820 3670 58848 4014
rect 58808 3664 58860 3670
rect 58808 3606 58860 3612
rect 58912 3602 58940 4134
rect 59452 4140 59504 4146
rect 59452 4082 59504 4088
rect 58716 3596 58768 3602
rect 58716 3538 58768 3544
rect 58900 3596 58952 3602
rect 58900 3538 58952 3544
rect 61016 3596 61068 3602
rect 61016 3538 61068 3544
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 58716 3392 58768 3398
rect 58716 3334 58768 3340
rect 57980 3120 58032 3126
rect 57980 3062 58032 3068
rect 56784 2916 56836 2922
rect 56784 2858 56836 2864
rect 57992 2650 58020 3062
rect 58728 3058 58756 3334
rect 58716 3052 58768 3058
rect 58716 2994 58768 3000
rect 59268 2916 59320 2922
rect 59268 2858 59320 2864
rect 57980 2644 58032 2650
rect 57980 2586 58032 2592
rect 58440 2576 58492 2582
rect 58440 2518 58492 2524
rect 57612 2440 57664 2446
rect 57612 2382 57664 2388
rect 57624 800 57652 2382
rect 58452 800 58480 2518
rect 59280 800 59308 2858
rect 60648 2848 60700 2854
rect 60648 2790 60700 2796
rect 60188 2508 60240 2514
rect 60188 2450 60240 2456
rect 60200 800 60228 2450
rect 60660 2378 60688 2790
rect 60648 2372 60700 2378
rect 60648 2314 60700 2320
rect 61028 800 61056 3538
rect 61936 3120 61988 3126
rect 61936 3062 61988 3068
rect 61948 800 61976 3062
rect 62764 2848 62816 2854
rect 62764 2790 62816 2796
rect 62776 800 62804 2790
rect 386 0 442 800
rect 1214 0 1270 800
rect 2042 0 2098 800
rect 2962 0 3018 800
rect 3790 0 3846 800
rect 4710 0 4766 800
rect 5538 0 5594 800
rect 6366 0 6422 800
rect 7286 0 7342 800
rect 8114 0 8170 800
rect 9034 0 9090 800
rect 9862 0 9918 800
rect 10782 0 10838 800
rect 11610 0 11666 800
rect 12438 0 12494 800
rect 13358 0 13414 800
rect 14186 0 14242 800
rect 15106 0 15162 800
rect 15934 0 15990 800
rect 16854 0 16910 800
rect 17682 0 17738 800
rect 18510 0 18566 800
rect 19430 0 19486 800
rect 20258 0 20314 800
rect 21178 0 21234 800
rect 22006 0 22062 800
rect 22926 0 22982 800
rect 23754 0 23810 800
rect 24582 0 24638 800
rect 25502 0 25558 800
rect 26330 0 26386 800
rect 27250 0 27306 800
rect 28078 0 28134 800
rect 28998 0 29054 800
rect 29826 0 29882 800
rect 30654 0 30710 800
rect 31574 0 31630 800
rect 32402 0 32458 800
rect 33322 0 33378 800
rect 34150 0 34206 800
rect 34978 0 35034 800
rect 35898 0 35954 800
rect 36726 0 36782 800
rect 37646 0 37702 800
rect 38474 0 38530 800
rect 39394 0 39450 800
rect 40222 0 40278 800
rect 41050 0 41106 800
rect 41970 0 42026 800
rect 42798 0 42854 800
rect 43718 0 43774 800
rect 44546 0 44602 800
rect 45466 0 45522 800
rect 46294 0 46350 800
rect 47122 0 47178 800
rect 48042 0 48098 800
rect 48870 0 48926 800
rect 49790 0 49846 800
rect 50618 0 50674 800
rect 51538 0 51594 800
rect 52366 0 52422 800
rect 53194 0 53250 800
rect 54114 0 54170 800
rect 54942 0 54998 800
rect 55862 0 55918 800
rect 56690 0 56746 800
rect 57610 0 57666 800
rect 58438 0 58494 800
rect 59266 0 59322 800
rect 60186 0 60242 800
rect 61014 0 61070 800
rect 61934 0 61990 800
rect 62762 0 62818 800
<< via2 >>
rect 3330 18536 3386 18592
rect 3054 16360 3110 16416
rect 4066 14184 4122 14240
rect 3514 12008 3570 12064
rect 2778 9832 2834 9888
rect 1858 6840 1914 6896
rect 2686 6196 2688 6216
rect 2688 6196 2740 6216
rect 2740 6196 2742 6216
rect 2686 6160 2742 6196
rect 2778 5480 2834 5536
rect 3054 7656 3110 7712
rect 1214 3712 1270 3768
rect 4066 3984 4122 4040
rect 3790 3440 3846 3496
rect 3422 1128 3478 1184
rect 4066 3304 4122 3360
rect 11137 17434 11193 17436
rect 11217 17434 11273 17436
rect 11297 17434 11353 17436
rect 11377 17434 11433 17436
rect 11137 17382 11163 17434
rect 11163 17382 11193 17434
rect 11217 17382 11227 17434
rect 11227 17382 11273 17434
rect 11297 17382 11343 17434
rect 11343 17382 11353 17434
rect 11377 17382 11407 17434
rect 11407 17382 11433 17434
rect 11137 17380 11193 17382
rect 11217 17380 11273 17382
rect 11297 17380 11353 17382
rect 11377 17380 11433 17382
rect 11137 16346 11193 16348
rect 11217 16346 11273 16348
rect 11297 16346 11353 16348
rect 11377 16346 11433 16348
rect 11137 16294 11163 16346
rect 11163 16294 11193 16346
rect 11217 16294 11227 16346
rect 11227 16294 11273 16346
rect 11297 16294 11343 16346
rect 11343 16294 11353 16346
rect 11377 16294 11407 16346
rect 11407 16294 11433 16346
rect 11137 16292 11193 16294
rect 11217 16292 11273 16294
rect 11297 16292 11353 16294
rect 11377 16292 11433 16294
rect 11137 15258 11193 15260
rect 11217 15258 11273 15260
rect 11297 15258 11353 15260
rect 11377 15258 11433 15260
rect 11137 15206 11163 15258
rect 11163 15206 11193 15258
rect 11217 15206 11227 15258
rect 11227 15206 11273 15258
rect 11297 15206 11343 15258
rect 11343 15206 11353 15258
rect 11377 15206 11407 15258
rect 11407 15206 11433 15258
rect 11137 15204 11193 15206
rect 11217 15204 11273 15206
rect 11297 15204 11353 15206
rect 11377 15204 11433 15206
rect 11137 14170 11193 14172
rect 11217 14170 11273 14172
rect 11297 14170 11353 14172
rect 11377 14170 11433 14172
rect 11137 14118 11163 14170
rect 11163 14118 11193 14170
rect 11217 14118 11227 14170
rect 11227 14118 11273 14170
rect 11297 14118 11343 14170
rect 11343 14118 11353 14170
rect 11377 14118 11407 14170
rect 11407 14118 11433 14170
rect 11137 14116 11193 14118
rect 11217 14116 11273 14118
rect 11297 14116 11353 14118
rect 11377 14116 11433 14118
rect 10966 13504 11022 13560
rect 5814 4684 5870 4720
rect 5814 4664 5816 4684
rect 5816 4664 5868 4684
rect 5868 4664 5870 4684
rect 4710 3032 4766 3088
rect 6366 3576 6422 3632
rect 5630 2896 5686 2952
rect 8758 10548 8760 10568
rect 8760 10548 8812 10568
rect 8812 10548 8814 10568
rect 8758 10512 8814 10548
rect 7838 5208 7894 5264
rect 9218 10512 9274 10568
rect 10782 13232 10838 13288
rect 9862 12280 9918 12336
rect 11137 13082 11193 13084
rect 11217 13082 11273 13084
rect 11297 13082 11353 13084
rect 11377 13082 11433 13084
rect 11137 13030 11163 13082
rect 11163 13030 11193 13082
rect 11217 13030 11227 13082
rect 11227 13030 11273 13082
rect 11297 13030 11343 13082
rect 11343 13030 11353 13082
rect 11377 13030 11407 13082
rect 11407 13030 11433 13082
rect 11137 13028 11193 13030
rect 11217 13028 11273 13030
rect 11297 13028 11353 13030
rect 11377 13028 11433 13030
rect 11137 11994 11193 11996
rect 11217 11994 11273 11996
rect 11297 11994 11353 11996
rect 11377 11994 11433 11996
rect 11137 11942 11163 11994
rect 11163 11942 11193 11994
rect 11217 11942 11227 11994
rect 11227 11942 11273 11994
rect 11297 11942 11343 11994
rect 11343 11942 11353 11994
rect 11377 11942 11407 11994
rect 11407 11942 11433 11994
rect 11137 11940 11193 11942
rect 11217 11940 11273 11942
rect 11297 11940 11353 11942
rect 11377 11940 11433 11942
rect 10782 11212 10838 11248
rect 10782 11192 10784 11212
rect 10784 11192 10836 11212
rect 10836 11192 10838 11212
rect 11242 11600 11298 11656
rect 11137 10906 11193 10908
rect 11217 10906 11273 10908
rect 11297 10906 11353 10908
rect 11377 10906 11433 10908
rect 11137 10854 11163 10906
rect 11163 10854 11193 10906
rect 11217 10854 11227 10906
rect 11227 10854 11273 10906
rect 11297 10854 11343 10906
rect 11343 10854 11353 10906
rect 11377 10854 11407 10906
rect 11407 10854 11433 10906
rect 11137 10852 11193 10854
rect 11217 10852 11273 10854
rect 11297 10852 11353 10854
rect 11377 10852 11433 10854
rect 11610 10784 11666 10840
rect 11137 9818 11193 9820
rect 11217 9818 11273 9820
rect 11297 9818 11353 9820
rect 11377 9818 11433 9820
rect 11137 9766 11163 9818
rect 11163 9766 11193 9818
rect 11217 9766 11227 9818
rect 11227 9766 11273 9818
rect 11297 9766 11343 9818
rect 11343 9766 11353 9818
rect 11377 9766 11407 9818
rect 11407 9766 11433 9818
rect 11137 9764 11193 9766
rect 11217 9764 11273 9766
rect 11297 9764 11353 9766
rect 11377 9764 11433 9766
rect 11137 8730 11193 8732
rect 11217 8730 11273 8732
rect 11297 8730 11353 8732
rect 11377 8730 11433 8732
rect 11137 8678 11163 8730
rect 11163 8678 11193 8730
rect 11217 8678 11227 8730
rect 11227 8678 11273 8730
rect 11297 8678 11343 8730
rect 11343 8678 11353 8730
rect 11377 8678 11407 8730
rect 11407 8678 11433 8730
rect 11137 8676 11193 8678
rect 11217 8676 11273 8678
rect 11297 8676 11353 8678
rect 11377 8676 11433 8678
rect 11137 7642 11193 7644
rect 11217 7642 11273 7644
rect 11297 7642 11353 7644
rect 11377 7642 11433 7644
rect 11137 7590 11163 7642
rect 11163 7590 11193 7642
rect 11217 7590 11227 7642
rect 11227 7590 11273 7642
rect 11297 7590 11343 7642
rect 11343 7590 11353 7642
rect 11377 7590 11407 7642
rect 11407 7590 11433 7642
rect 11137 7588 11193 7590
rect 11217 7588 11273 7590
rect 11297 7588 11353 7590
rect 11377 7588 11433 7590
rect 11137 6554 11193 6556
rect 11217 6554 11273 6556
rect 11297 6554 11353 6556
rect 11377 6554 11433 6556
rect 11137 6502 11163 6554
rect 11163 6502 11193 6554
rect 11217 6502 11227 6554
rect 11227 6502 11273 6554
rect 11297 6502 11343 6554
rect 11343 6502 11353 6554
rect 11377 6502 11407 6554
rect 11407 6502 11433 6554
rect 11137 6500 11193 6502
rect 11217 6500 11273 6502
rect 11297 6500 11353 6502
rect 11377 6500 11433 6502
rect 12346 11772 12348 11792
rect 12348 11772 12400 11792
rect 12400 11772 12402 11792
rect 12346 11736 12402 11772
rect 12346 9036 12402 9072
rect 12346 9016 12348 9036
rect 12348 9016 12400 9036
rect 12400 9016 12402 9036
rect 11137 5466 11193 5468
rect 11217 5466 11273 5468
rect 11297 5466 11353 5468
rect 11377 5466 11433 5468
rect 11137 5414 11163 5466
rect 11163 5414 11193 5466
rect 11217 5414 11227 5466
rect 11227 5414 11273 5466
rect 11297 5414 11343 5466
rect 11343 5414 11353 5466
rect 11377 5414 11407 5466
rect 11407 5414 11433 5466
rect 11137 5412 11193 5414
rect 11217 5412 11273 5414
rect 11297 5412 11353 5414
rect 11377 5412 11433 5414
rect 10966 5072 11022 5128
rect 12898 11872 12954 11928
rect 13266 11736 13322 11792
rect 13174 11464 13230 11520
rect 12622 7948 12678 7984
rect 12622 7928 12624 7948
rect 12624 7928 12676 7948
rect 12676 7928 12678 7948
rect 12162 4528 12218 4584
rect 11137 4378 11193 4380
rect 11217 4378 11273 4380
rect 11297 4378 11353 4380
rect 11377 4378 11433 4380
rect 11137 4326 11163 4378
rect 11163 4326 11193 4378
rect 11217 4326 11227 4378
rect 11227 4326 11273 4378
rect 11297 4326 11343 4378
rect 11343 4326 11353 4378
rect 11377 4326 11407 4378
rect 11407 4326 11433 4378
rect 11137 4324 11193 4326
rect 11217 4324 11273 4326
rect 11297 4324 11353 4326
rect 11377 4324 11433 4326
rect 9954 4120 10010 4176
rect 10690 4120 10746 4176
rect 9770 3712 9826 3768
rect 11137 3290 11193 3292
rect 11217 3290 11273 3292
rect 11297 3290 11353 3292
rect 11377 3290 11433 3292
rect 11137 3238 11163 3290
rect 11163 3238 11193 3290
rect 11217 3238 11227 3290
rect 11227 3238 11273 3290
rect 11297 3238 11343 3290
rect 11343 3238 11353 3290
rect 11377 3238 11407 3290
rect 11407 3238 11433 3290
rect 11137 3236 11193 3238
rect 11217 3236 11273 3238
rect 11297 3236 11353 3238
rect 11377 3236 11433 3238
rect 11137 2202 11193 2204
rect 11217 2202 11273 2204
rect 11297 2202 11353 2204
rect 11377 2202 11433 2204
rect 11137 2150 11163 2202
rect 11163 2150 11193 2202
rect 11217 2150 11227 2202
rect 11227 2150 11273 2202
rect 11297 2150 11343 2202
rect 11343 2150 11353 2202
rect 11377 2150 11407 2202
rect 11407 2150 11433 2202
rect 11137 2148 11193 2150
rect 11217 2148 11273 2150
rect 11297 2148 11353 2150
rect 11377 2148 11433 2150
rect 12806 4664 12862 4720
rect 13358 11600 13414 11656
rect 16578 13504 16634 13560
rect 15290 13232 15346 13288
rect 14554 11192 14610 11248
rect 13450 5208 13506 5264
rect 14738 3304 14794 3360
rect 16394 11872 16450 11928
rect 17774 12300 17830 12336
rect 17774 12280 17776 12300
rect 17776 12280 17828 12300
rect 17828 12280 17830 12300
rect 21318 16890 21374 16892
rect 21398 16890 21454 16892
rect 21478 16890 21534 16892
rect 21558 16890 21614 16892
rect 21318 16838 21344 16890
rect 21344 16838 21374 16890
rect 21398 16838 21408 16890
rect 21408 16838 21454 16890
rect 21478 16838 21524 16890
rect 21524 16838 21534 16890
rect 21558 16838 21588 16890
rect 21588 16838 21614 16890
rect 21318 16836 21374 16838
rect 21398 16836 21454 16838
rect 21478 16836 21534 16838
rect 21558 16836 21614 16838
rect 19430 13368 19486 13424
rect 19062 13232 19118 13288
rect 18878 11872 18934 11928
rect 18786 11464 18842 11520
rect 19338 10004 19340 10024
rect 19340 10004 19392 10024
rect 19392 10004 19394 10024
rect 19338 9968 19394 10004
rect 15290 3848 15346 3904
rect 17958 9016 18014 9072
rect 17774 8916 17776 8936
rect 17776 8916 17828 8936
rect 17828 8916 17830 8936
rect 17774 8880 17830 8916
rect 16578 2624 16634 2680
rect 17222 3304 17278 3360
rect 16762 2760 16818 2816
rect 17866 7964 17868 7984
rect 17868 7964 17920 7984
rect 17920 7964 17922 7984
rect 17866 7928 17922 7964
rect 21318 15802 21374 15804
rect 21398 15802 21454 15804
rect 21478 15802 21534 15804
rect 21558 15802 21614 15804
rect 21318 15750 21344 15802
rect 21344 15750 21374 15802
rect 21398 15750 21408 15802
rect 21408 15750 21454 15802
rect 21478 15750 21524 15802
rect 21524 15750 21534 15802
rect 21558 15750 21588 15802
rect 21588 15750 21614 15802
rect 21318 15748 21374 15750
rect 21398 15748 21454 15750
rect 21478 15748 21534 15750
rect 21558 15748 21614 15750
rect 21318 14714 21374 14716
rect 21398 14714 21454 14716
rect 21478 14714 21534 14716
rect 21558 14714 21614 14716
rect 21318 14662 21344 14714
rect 21344 14662 21374 14714
rect 21398 14662 21408 14714
rect 21408 14662 21454 14714
rect 21478 14662 21524 14714
rect 21524 14662 21534 14714
rect 21558 14662 21588 14714
rect 21588 14662 21614 14714
rect 21318 14660 21374 14662
rect 21398 14660 21454 14662
rect 21478 14660 21534 14662
rect 21558 14660 21614 14662
rect 19614 9596 19616 9616
rect 19616 9596 19668 9616
rect 19668 9596 19670 9616
rect 19614 9560 19670 9596
rect 20350 13096 20406 13152
rect 20442 12960 20498 13016
rect 21318 13626 21374 13628
rect 21398 13626 21454 13628
rect 21478 13626 21534 13628
rect 21558 13626 21614 13628
rect 21318 13574 21344 13626
rect 21344 13574 21374 13626
rect 21398 13574 21408 13626
rect 21408 13574 21454 13626
rect 21478 13574 21524 13626
rect 21524 13574 21534 13626
rect 21558 13574 21588 13626
rect 21588 13574 21614 13626
rect 21318 13572 21374 13574
rect 21398 13572 21454 13574
rect 21478 13572 21534 13574
rect 21558 13572 21614 13574
rect 20810 11756 20866 11792
rect 20810 11736 20812 11756
rect 20812 11736 20864 11756
rect 20864 11736 20866 11756
rect 21086 11192 21142 11248
rect 20902 11092 20904 11112
rect 20904 11092 20956 11112
rect 20956 11092 20958 11112
rect 20902 11056 20958 11092
rect 20902 10804 20958 10840
rect 20902 10784 20904 10804
rect 20904 10784 20956 10804
rect 20956 10784 20958 10804
rect 20994 9968 21050 10024
rect 20810 9696 20866 9752
rect 21318 12538 21374 12540
rect 21398 12538 21454 12540
rect 21478 12538 21534 12540
rect 21558 12538 21614 12540
rect 21318 12486 21344 12538
rect 21344 12486 21374 12538
rect 21398 12486 21408 12538
rect 21408 12486 21454 12538
rect 21478 12486 21524 12538
rect 21524 12486 21534 12538
rect 21558 12486 21588 12538
rect 21588 12486 21614 12538
rect 21318 12484 21374 12486
rect 21398 12484 21454 12486
rect 21478 12484 21534 12486
rect 21558 12484 21614 12486
rect 21318 11450 21374 11452
rect 21398 11450 21454 11452
rect 21478 11450 21534 11452
rect 21558 11450 21614 11452
rect 21318 11398 21344 11450
rect 21344 11398 21374 11450
rect 21398 11398 21408 11450
rect 21408 11398 21454 11450
rect 21478 11398 21524 11450
rect 21524 11398 21534 11450
rect 21558 11398 21588 11450
rect 21588 11398 21614 11450
rect 21318 11396 21374 11398
rect 21398 11396 21454 11398
rect 21478 11396 21534 11398
rect 21558 11396 21614 11398
rect 22650 12824 22706 12880
rect 21318 10362 21374 10364
rect 21398 10362 21454 10364
rect 21478 10362 21534 10364
rect 21558 10362 21614 10364
rect 21318 10310 21344 10362
rect 21344 10310 21374 10362
rect 21398 10310 21408 10362
rect 21408 10310 21454 10362
rect 21478 10310 21524 10362
rect 21524 10310 21534 10362
rect 21558 10310 21588 10362
rect 21588 10310 21614 10362
rect 21318 10308 21374 10310
rect 21398 10308 21454 10310
rect 21478 10308 21534 10310
rect 21558 10308 21614 10310
rect 20258 9016 20314 9072
rect 18234 4256 18290 4312
rect 18786 4528 18842 4584
rect 18970 4528 19026 4584
rect 19246 4256 19302 4312
rect 19338 4120 19394 4176
rect 18694 2760 18750 2816
rect 18786 2624 18842 2680
rect 19154 3848 19210 3904
rect 20166 8492 20222 8528
rect 20166 8472 20168 8492
rect 20168 8472 20220 8492
rect 20220 8472 20222 8492
rect 21318 9274 21374 9276
rect 21398 9274 21454 9276
rect 21478 9274 21534 9276
rect 21558 9274 21614 9276
rect 21318 9222 21344 9274
rect 21344 9222 21374 9274
rect 21398 9222 21408 9274
rect 21408 9222 21454 9274
rect 21478 9222 21524 9274
rect 21524 9222 21534 9274
rect 21558 9222 21588 9274
rect 21588 9222 21614 9274
rect 21318 9220 21374 9222
rect 21398 9220 21454 9222
rect 21478 9220 21534 9222
rect 21558 9220 21614 9222
rect 21546 9036 21602 9072
rect 21546 9016 21548 9036
rect 21548 9016 21600 9036
rect 21600 9016 21602 9036
rect 20902 8880 20958 8936
rect 20718 8608 20774 8664
rect 20442 7792 20498 7848
rect 20074 6432 20130 6488
rect 20350 6296 20406 6352
rect 21318 8186 21374 8188
rect 21398 8186 21454 8188
rect 21478 8186 21534 8188
rect 21558 8186 21614 8188
rect 21318 8134 21344 8186
rect 21344 8134 21374 8186
rect 21398 8134 21408 8186
rect 21408 8134 21454 8186
rect 21478 8134 21524 8186
rect 21524 8134 21534 8186
rect 21558 8134 21588 8186
rect 21588 8134 21614 8186
rect 21318 8132 21374 8134
rect 21398 8132 21454 8134
rect 21478 8132 21534 8134
rect 21558 8132 21614 8134
rect 20994 6704 21050 6760
rect 20534 3984 20590 4040
rect 21318 7098 21374 7100
rect 21398 7098 21454 7100
rect 21478 7098 21534 7100
rect 21558 7098 21614 7100
rect 21318 7046 21344 7098
rect 21344 7046 21374 7098
rect 21398 7046 21408 7098
rect 21408 7046 21454 7098
rect 21478 7046 21524 7098
rect 21524 7046 21534 7098
rect 21558 7046 21588 7098
rect 21588 7046 21614 7098
rect 21318 7044 21374 7046
rect 21398 7044 21454 7046
rect 21478 7044 21534 7046
rect 21558 7044 21614 7046
rect 21822 8356 21878 8392
rect 21822 8336 21824 8356
rect 21824 8336 21876 8356
rect 21876 8336 21878 8356
rect 22006 8472 22062 8528
rect 22558 8608 22614 8664
rect 21730 6160 21786 6216
rect 21318 6010 21374 6012
rect 21398 6010 21454 6012
rect 21478 6010 21534 6012
rect 21558 6010 21614 6012
rect 21318 5958 21344 6010
rect 21344 5958 21374 6010
rect 21398 5958 21408 6010
rect 21408 5958 21454 6010
rect 21478 5958 21524 6010
rect 21524 5958 21534 6010
rect 21558 5958 21588 6010
rect 21588 5958 21614 6010
rect 21318 5956 21374 5958
rect 21398 5956 21454 5958
rect 21478 5956 21534 5958
rect 21558 5956 21614 5958
rect 21178 5480 21234 5536
rect 21318 4922 21374 4924
rect 21398 4922 21454 4924
rect 21478 4922 21534 4924
rect 21558 4922 21614 4924
rect 21318 4870 21344 4922
rect 21344 4870 21374 4922
rect 21398 4870 21408 4922
rect 21408 4870 21454 4922
rect 21478 4870 21524 4922
rect 21524 4870 21534 4922
rect 21558 4870 21588 4922
rect 21588 4870 21614 4922
rect 21318 4868 21374 4870
rect 21398 4868 21454 4870
rect 21478 4868 21534 4870
rect 21558 4868 21614 4870
rect 21318 3834 21374 3836
rect 21398 3834 21454 3836
rect 21478 3834 21534 3836
rect 21558 3834 21614 3836
rect 21318 3782 21344 3834
rect 21344 3782 21374 3834
rect 21398 3782 21408 3834
rect 21408 3782 21454 3834
rect 21478 3782 21524 3834
rect 21524 3782 21534 3834
rect 21558 3782 21588 3834
rect 21588 3782 21614 3834
rect 21318 3780 21374 3782
rect 21398 3780 21454 3782
rect 21478 3780 21534 3782
rect 21558 3780 21614 3782
rect 22006 3304 22062 3360
rect 21318 2746 21374 2748
rect 21398 2746 21454 2748
rect 21478 2746 21534 2748
rect 21558 2746 21614 2748
rect 21318 2694 21344 2746
rect 21344 2694 21374 2746
rect 21398 2694 21408 2746
rect 21408 2694 21454 2746
rect 21478 2694 21524 2746
rect 21524 2694 21534 2746
rect 21558 2694 21588 2746
rect 21588 2694 21614 2746
rect 21318 2692 21374 2694
rect 21398 2692 21454 2694
rect 21478 2692 21534 2694
rect 21558 2692 21614 2694
rect 23018 13388 23074 13424
rect 23018 13368 23020 13388
rect 23020 13368 23072 13388
rect 23072 13368 23074 13388
rect 23754 11772 23756 11792
rect 23756 11772 23808 11792
rect 23808 11772 23810 11792
rect 23754 11736 23810 11772
rect 23754 9596 23756 9616
rect 23756 9596 23808 9616
rect 23808 9596 23810 9616
rect 23754 9560 23810 9596
rect 31500 17434 31556 17436
rect 31580 17434 31636 17436
rect 31660 17434 31716 17436
rect 31740 17434 31796 17436
rect 31500 17382 31526 17434
rect 31526 17382 31556 17434
rect 31580 17382 31590 17434
rect 31590 17382 31636 17434
rect 31660 17382 31706 17434
rect 31706 17382 31716 17434
rect 31740 17382 31770 17434
rect 31770 17382 31796 17434
rect 31500 17380 31556 17382
rect 31580 17380 31636 17382
rect 31660 17380 31716 17382
rect 31740 17380 31796 17382
rect 31500 16346 31556 16348
rect 31580 16346 31636 16348
rect 31660 16346 31716 16348
rect 31740 16346 31796 16348
rect 31500 16294 31526 16346
rect 31526 16294 31556 16346
rect 31580 16294 31590 16346
rect 31590 16294 31636 16346
rect 31660 16294 31706 16346
rect 31706 16294 31716 16346
rect 31740 16294 31770 16346
rect 31770 16294 31796 16346
rect 31500 16292 31556 16294
rect 31580 16292 31636 16294
rect 31660 16292 31716 16294
rect 31740 16292 31796 16294
rect 24950 11056 25006 11112
rect 27066 13096 27122 13152
rect 26882 12960 26938 13016
rect 26330 12552 26386 12608
rect 27710 12824 27766 12880
rect 27894 12588 27896 12608
rect 27896 12588 27948 12608
rect 27948 12588 27950 12608
rect 27894 12552 27950 12588
rect 25226 9560 25282 9616
rect 27802 11192 27858 11248
rect 22650 7792 22706 7848
rect 22926 3984 22982 4040
rect 22558 3032 22614 3088
rect 22374 2896 22430 2952
rect 24030 5208 24086 5264
rect 23938 4120 23994 4176
rect 24582 3712 24638 3768
rect 23754 3168 23810 3224
rect 24122 2624 24178 2680
rect 27158 8336 27214 8392
rect 25502 5108 25504 5128
rect 25504 5108 25556 5128
rect 25556 5108 25558 5128
rect 25502 5072 25558 5108
rect 27158 5908 27214 5944
rect 27710 9016 27766 9072
rect 28078 6976 28134 7032
rect 27158 5888 27160 5908
rect 27160 5888 27212 5908
rect 27212 5888 27214 5908
rect 26790 3848 26846 3904
rect 26790 3304 26846 3360
rect 26330 2896 26386 2952
rect 26974 3576 27030 3632
rect 26974 2760 27030 2816
rect 28262 5480 28318 5536
rect 28630 10512 28686 10568
rect 28538 6432 28594 6488
rect 29366 12708 29422 12744
rect 29366 12688 29368 12708
rect 29368 12688 29420 12708
rect 29420 12688 29422 12708
rect 30010 12436 30066 12472
rect 30010 12416 30012 12436
rect 30012 12416 30064 12436
rect 30064 12416 30066 12436
rect 28814 5516 28816 5536
rect 28816 5516 28868 5536
rect 28868 5516 28870 5536
rect 28814 5480 28870 5516
rect 27342 3576 27398 3632
rect 29366 5480 29422 5536
rect 31500 15258 31556 15260
rect 31580 15258 31636 15260
rect 31660 15258 31716 15260
rect 31740 15258 31796 15260
rect 31500 15206 31526 15258
rect 31526 15206 31556 15258
rect 31580 15206 31590 15258
rect 31590 15206 31636 15258
rect 31660 15206 31706 15258
rect 31706 15206 31716 15258
rect 31740 15206 31770 15258
rect 31770 15206 31796 15258
rect 31500 15204 31556 15206
rect 31580 15204 31636 15206
rect 31660 15204 31716 15206
rect 31740 15204 31796 15206
rect 31500 14170 31556 14172
rect 31580 14170 31636 14172
rect 31660 14170 31716 14172
rect 31740 14170 31796 14172
rect 31500 14118 31526 14170
rect 31526 14118 31556 14170
rect 31580 14118 31590 14170
rect 31590 14118 31636 14170
rect 31660 14118 31706 14170
rect 31706 14118 31716 14170
rect 31740 14118 31770 14170
rect 31770 14118 31796 14170
rect 31500 14116 31556 14118
rect 31580 14116 31636 14118
rect 31660 14116 31716 14118
rect 31740 14116 31796 14118
rect 30470 12180 30472 12200
rect 30472 12180 30524 12200
rect 30524 12180 30526 12200
rect 30470 12144 30526 12180
rect 31500 13082 31556 13084
rect 31580 13082 31636 13084
rect 31660 13082 31716 13084
rect 31740 13082 31796 13084
rect 31500 13030 31526 13082
rect 31526 13030 31556 13082
rect 31580 13030 31590 13082
rect 31590 13030 31636 13082
rect 31660 13030 31706 13082
rect 31706 13030 31716 13082
rect 31740 13030 31770 13082
rect 31770 13030 31796 13082
rect 31500 13028 31556 13030
rect 31580 13028 31636 13030
rect 31660 13028 31716 13030
rect 31740 13028 31796 13030
rect 31206 12180 31208 12200
rect 31208 12180 31260 12200
rect 31260 12180 31262 12200
rect 31206 12144 31262 12180
rect 31500 11994 31556 11996
rect 31580 11994 31636 11996
rect 31660 11994 31716 11996
rect 31740 11994 31796 11996
rect 31500 11942 31526 11994
rect 31526 11942 31556 11994
rect 31580 11942 31590 11994
rect 31590 11942 31636 11994
rect 31660 11942 31706 11994
rect 31706 11942 31716 11994
rect 31740 11942 31770 11994
rect 31770 11942 31796 11994
rect 31500 11940 31556 11942
rect 31580 11940 31636 11942
rect 31660 11940 31716 11942
rect 31740 11940 31796 11942
rect 33874 12824 33930 12880
rect 34242 12688 34298 12744
rect 30194 7112 30250 7168
rect 30286 6024 30342 6080
rect 30194 4800 30250 4856
rect 29826 3032 29882 3088
rect 30562 5616 30618 5672
rect 30930 5772 30986 5808
rect 30930 5752 30932 5772
rect 30932 5752 30984 5772
rect 30984 5752 30986 5772
rect 31500 10906 31556 10908
rect 31580 10906 31636 10908
rect 31660 10906 31716 10908
rect 31740 10906 31796 10908
rect 31500 10854 31526 10906
rect 31526 10854 31556 10906
rect 31580 10854 31590 10906
rect 31590 10854 31636 10906
rect 31660 10854 31706 10906
rect 31706 10854 31716 10906
rect 31740 10854 31770 10906
rect 31770 10854 31796 10906
rect 31500 10852 31556 10854
rect 31580 10852 31636 10854
rect 31660 10852 31716 10854
rect 31740 10852 31796 10854
rect 31500 9818 31556 9820
rect 31580 9818 31636 9820
rect 31660 9818 31716 9820
rect 31740 9818 31796 9820
rect 31500 9766 31526 9818
rect 31526 9766 31556 9818
rect 31580 9766 31590 9818
rect 31590 9766 31636 9818
rect 31660 9766 31706 9818
rect 31706 9766 31716 9818
rect 31740 9766 31770 9818
rect 31770 9766 31796 9818
rect 31500 9764 31556 9766
rect 31580 9764 31636 9766
rect 31660 9764 31716 9766
rect 31740 9764 31796 9766
rect 31298 9696 31354 9752
rect 31500 8730 31556 8732
rect 31580 8730 31636 8732
rect 31660 8730 31716 8732
rect 31740 8730 31796 8732
rect 31500 8678 31526 8730
rect 31526 8678 31556 8730
rect 31580 8678 31590 8730
rect 31590 8678 31636 8730
rect 31660 8678 31706 8730
rect 31706 8678 31716 8730
rect 31740 8678 31770 8730
rect 31770 8678 31796 8730
rect 31500 8676 31556 8678
rect 31580 8676 31636 8678
rect 31660 8676 31716 8678
rect 31740 8676 31796 8678
rect 31850 8492 31906 8528
rect 31850 8472 31852 8492
rect 31852 8472 31904 8492
rect 31904 8472 31906 8492
rect 32126 8472 32182 8528
rect 31500 7642 31556 7644
rect 31580 7642 31636 7644
rect 31660 7642 31716 7644
rect 31740 7642 31796 7644
rect 31500 7590 31526 7642
rect 31526 7590 31556 7642
rect 31580 7590 31590 7642
rect 31590 7590 31636 7642
rect 31660 7590 31706 7642
rect 31706 7590 31716 7642
rect 31740 7590 31770 7642
rect 31770 7590 31796 7642
rect 31500 7588 31556 7590
rect 31580 7588 31636 7590
rect 31660 7588 31716 7590
rect 31740 7588 31796 7590
rect 31206 6196 31208 6216
rect 31208 6196 31260 6216
rect 31260 6196 31262 6216
rect 31206 6160 31262 6196
rect 31022 4528 31078 4584
rect 30654 3984 30710 4040
rect 30378 2624 30434 2680
rect 31298 5908 31354 5944
rect 31298 5888 31300 5908
rect 31300 5888 31352 5908
rect 31352 5888 31354 5908
rect 32034 6976 32090 7032
rect 32218 7928 32274 7984
rect 31500 6554 31556 6556
rect 31580 6554 31636 6556
rect 31660 6554 31716 6556
rect 31740 6554 31796 6556
rect 31500 6502 31526 6554
rect 31526 6502 31556 6554
rect 31580 6502 31590 6554
rect 31590 6502 31636 6554
rect 31660 6502 31706 6554
rect 31706 6502 31716 6554
rect 31740 6502 31770 6554
rect 31770 6502 31796 6554
rect 31500 6500 31556 6502
rect 31580 6500 31636 6502
rect 31660 6500 31716 6502
rect 31740 6500 31796 6502
rect 31758 6024 31814 6080
rect 31850 5636 31906 5672
rect 31850 5616 31852 5636
rect 31852 5616 31904 5636
rect 31904 5616 31906 5636
rect 31500 5466 31556 5468
rect 31580 5466 31636 5468
rect 31660 5466 31716 5468
rect 31740 5466 31796 5468
rect 31500 5414 31526 5466
rect 31526 5414 31556 5466
rect 31580 5414 31590 5466
rect 31590 5414 31636 5466
rect 31660 5414 31706 5466
rect 31706 5414 31716 5466
rect 31740 5414 31770 5466
rect 31770 5414 31796 5466
rect 31500 5412 31556 5414
rect 31580 5412 31636 5414
rect 31660 5412 31716 5414
rect 31740 5412 31796 5414
rect 31500 4378 31556 4380
rect 31580 4378 31636 4380
rect 31660 4378 31716 4380
rect 31740 4378 31796 4380
rect 31500 4326 31526 4378
rect 31526 4326 31556 4378
rect 31580 4326 31590 4378
rect 31590 4326 31636 4378
rect 31660 4326 31706 4378
rect 31706 4326 31716 4378
rect 31740 4326 31770 4378
rect 31770 4326 31796 4378
rect 31500 4324 31556 4326
rect 31580 4324 31636 4326
rect 31660 4324 31716 4326
rect 31740 4324 31796 4326
rect 31666 3712 31722 3768
rect 31850 3712 31906 3768
rect 31942 3304 31998 3360
rect 31500 3290 31556 3292
rect 31580 3290 31636 3292
rect 31660 3290 31716 3292
rect 31740 3290 31796 3292
rect 31500 3238 31526 3290
rect 31526 3238 31556 3290
rect 31580 3238 31590 3290
rect 31590 3238 31636 3290
rect 31660 3238 31706 3290
rect 31706 3238 31716 3290
rect 31740 3238 31770 3290
rect 31770 3238 31796 3290
rect 31500 3236 31556 3238
rect 31580 3236 31636 3238
rect 31660 3236 31716 3238
rect 31740 3236 31796 3238
rect 31298 3168 31354 3224
rect 32402 5788 32404 5808
rect 32404 5788 32456 5808
rect 32456 5788 32458 5808
rect 32402 5752 32458 5788
rect 32954 7928 33010 7984
rect 32862 7248 32918 7304
rect 32770 6704 32826 6760
rect 32586 6160 32642 6216
rect 32494 4800 32550 4856
rect 32310 2760 32366 2816
rect 31500 2202 31556 2204
rect 31580 2202 31636 2204
rect 31660 2202 31716 2204
rect 31740 2202 31796 2204
rect 31500 2150 31526 2202
rect 31526 2150 31556 2202
rect 31580 2150 31590 2202
rect 31590 2150 31636 2202
rect 31660 2150 31706 2202
rect 31706 2150 31716 2202
rect 31740 2150 31770 2202
rect 31770 2150 31796 2202
rect 31500 2148 31556 2150
rect 31580 2148 31636 2150
rect 31660 2148 31716 2150
rect 31740 2148 31796 2150
rect 36082 12824 36138 12880
rect 32954 4120 33010 4176
rect 37370 12416 37426 12472
rect 35714 6976 35770 7032
rect 35990 7112 36046 7168
rect 34242 3168 34298 3224
rect 33966 2624 34022 2680
rect 34702 3576 34758 3632
rect 34518 3304 34574 3360
rect 34702 3304 34758 3360
rect 34518 2760 34574 2816
rect 41681 16890 41737 16892
rect 41761 16890 41817 16892
rect 41841 16890 41897 16892
rect 41921 16890 41977 16892
rect 41681 16838 41707 16890
rect 41707 16838 41737 16890
rect 41761 16838 41771 16890
rect 41771 16838 41817 16890
rect 41841 16838 41887 16890
rect 41887 16838 41897 16890
rect 41921 16838 41951 16890
rect 41951 16838 41977 16890
rect 41681 16836 41737 16838
rect 41761 16836 41817 16838
rect 41841 16836 41897 16838
rect 41921 16836 41977 16838
rect 41681 15802 41737 15804
rect 41761 15802 41817 15804
rect 41841 15802 41897 15804
rect 41921 15802 41977 15804
rect 41681 15750 41707 15802
rect 41707 15750 41737 15802
rect 41761 15750 41771 15802
rect 41771 15750 41817 15802
rect 41841 15750 41887 15802
rect 41887 15750 41897 15802
rect 41921 15750 41951 15802
rect 41951 15750 41977 15802
rect 41681 15748 41737 15750
rect 41761 15748 41817 15750
rect 41841 15748 41897 15750
rect 41921 15748 41977 15750
rect 37278 9580 37334 9616
rect 37278 9560 37280 9580
rect 37280 9560 37332 9580
rect 37332 9560 37334 9580
rect 35346 4548 35402 4584
rect 35346 4528 35348 4548
rect 35348 4528 35400 4548
rect 35400 4528 35402 4548
rect 34978 3576 35034 3632
rect 35530 3476 35532 3496
rect 35532 3476 35584 3496
rect 35584 3476 35586 3496
rect 35530 3440 35586 3476
rect 36266 3712 36322 3768
rect 36174 2624 36230 2680
rect 37278 6704 37334 6760
rect 36818 3848 36874 3904
rect 39670 11872 39726 11928
rect 38566 7148 38568 7168
rect 38568 7148 38620 7168
rect 38620 7148 38622 7168
rect 38566 7112 38622 7148
rect 38750 7112 38806 7168
rect 36542 2760 36598 2816
rect 39026 3440 39082 3496
rect 41681 14714 41737 14716
rect 41761 14714 41817 14716
rect 41841 14714 41897 14716
rect 41921 14714 41977 14716
rect 41681 14662 41707 14714
rect 41707 14662 41737 14714
rect 41761 14662 41771 14714
rect 41771 14662 41817 14714
rect 41841 14662 41887 14714
rect 41887 14662 41897 14714
rect 41921 14662 41951 14714
rect 41951 14662 41977 14714
rect 41681 14660 41737 14662
rect 41761 14660 41817 14662
rect 41841 14660 41897 14662
rect 41921 14660 41977 14662
rect 41681 13626 41737 13628
rect 41761 13626 41817 13628
rect 41841 13626 41897 13628
rect 41921 13626 41977 13628
rect 41681 13574 41707 13626
rect 41707 13574 41737 13626
rect 41761 13574 41771 13626
rect 41771 13574 41817 13626
rect 41841 13574 41887 13626
rect 41887 13574 41897 13626
rect 41921 13574 41951 13626
rect 41951 13574 41977 13626
rect 41681 13572 41737 13574
rect 41761 13572 41817 13574
rect 41841 13572 41897 13574
rect 41921 13572 41977 13574
rect 41234 11600 41290 11656
rect 41418 9560 41474 9616
rect 41681 12538 41737 12540
rect 41761 12538 41817 12540
rect 41841 12538 41897 12540
rect 41921 12538 41977 12540
rect 41681 12486 41707 12538
rect 41707 12486 41737 12538
rect 41761 12486 41771 12538
rect 41771 12486 41817 12538
rect 41841 12486 41887 12538
rect 41887 12486 41897 12538
rect 41921 12486 41951 12538
rect 41951 12486 41977 12538
rect 41681 12484 41737 12486
rect 41761 12484 41817 12486
rect 41841 12484 41897 12486
rect 41921 12484 41977 12486
rect 41681 11450 41737 11452
rect 41761 11450 41817 11452
rect 41841 11450 41897 11452
rect 41921 11450 41977 11452
rect 41681 11398 41707 11450
rect 41707 11398 41737 11450
rect 41761 11398 41771 11450
rect 41771 11398 41817 11450
rect 41841 11398 41887 11450
rect 41887 11398 41897 11450
rect 41921 11398 41951 11450
rect 41951 11398 41977 11450
rect 41681 11396 41737 11398
rect 41761 11396 41817 11398
rect 41841 11396 41897 11398
rect 41921 11396 41977 11398
rect 41681 10362 41737 10364
rect 41761 10362 41817 10364
rect 41841 10362 41897 10364
rect 41921 10362 41977 10364
rect 41681 10310 41707 10362
rect 41707 10310 41737 10362
rect 41761 10310 41771 10362
rect 41771 10310 41817 10362
rect 41841 10310 41887 10362
rect 41887 10310 41897 10362
rect 41921 10310 41951 10362
rect 41951 10310 41977 10362
rect 41681 10308 41737 10310
rect 41761 10308 41817 10310
rect 41841 10308 41897 10310
rect 41921 10308 41977 10310
rect 41681 9274 41737 9276
rect 41761 9274 41817 9276
rect 41841 9274 41897 9276
rect 41921 9274 41977 9276
rect 41681 9222 41707 9274
rect 41707 9222 41737 9274
rect 41761 9222 41771 9274
rect 41771 9222 41817 9274
rect 41841 9222 41887 9274
rect 41887 9222 41897 9274
rect 41921 9222 41951 9274
rect 41951 9222 41977 9274
rect 41681 9220 41737 9222
rect 41761 9220 41817 9222
rect 41841 9220 41897 9222
rect 41921 9220 41977 9222
rect 40958 8336 41014 8392
rect 41234 8336 41290 8392
rect 40866 7384 40922 7440
rect 42154 8608 42210 8664
rect 42154 8200 42210 8256
rect 41681 8186 41737 8188
rect 41761 8186 41817 8188
rect 41841 8186 41897 8188
rect 41921 8186 41977 8188
rect 41681 8134 41707 8186
rect 41707 8134 41737 8186
rect 41761 8134 41771 8186
rect 41771 8134 41817 8186
rect 41841 8134 41887 8186
rect 41887 8134 41897 8186
rect 41921 8134 41951 8186
rect 41951 8134 41977 8186
rect 41681 8132 41737 8134
rect 41761 8132 41817 8134
rect 41841 8132 41897 8134
rect 41921 8132 41977 8134
rect 41234 6976 41290 7032
rect 41681 7098 41737 7100
rect 41761 7098 41817 7100
rect 41841 7098 41897 7100
rect 41921 7098 41977 7100
rect 41681 7046 41707 7098
rect 41707 7046 41737 7098
rect 41761 7046 41771 7098
rect 41771 7046 41817 7098
rect 41841 7046 41887 7098
rect 41887 7046 41897 7098
rect 41921 7046 41951 7098
rect 41951 7046 41977 7098
rect 41681 7044 41737 7046
rect 41761 7044 41817 7046
rect 41841 7044 41897 7046
rect 41921 7044 41977 7046
rect 41694 6432 41750 6488
rect 42154 6296 42210 6352
rect 41681 6010 41737 6012
rect 41761 6010 41817 6012
rect 41841 6010 41897 6012
rect 41921 6010 41977 6012
rect 41681 5958 41707 6010
rect 41707 5958 41737 6010
rect 41761 5958 41771 6010
rect 41771 5958 41817 6010
rect 41841 5958 41887 6010
rect 41887 5958 41897 6010
rect 41921 5958 41951 6010
rect 41951 5958 41977 6010
rect 41681 5956 41737 5958
rect 41761 5956 41817 5958
rect 41841 5956 41897 5958
rect 41921 5956 41977 5958
rect 41418 5208 41474 5264
rect 41681 4922 41737 4924
rect 41761 4922 41817 4924
rect 41841 4922 41897 4924
rect 41921 4922 41977 4924
rect 41681 4870 41707 4922
rect 41707 4870 41737 4922
rect 41761 4870 41771 4922
rect 41771 4870 41817 4922
rect 41841 4870 41887 4922
rect 41887 4870 41897 4922
rect 41921 4870 41951 4922
rect 41951 4870 41977 4922
rect 41681 4868 41737 4870
rect 41761 4868 41817 4870
rect 41841 4868 41897 4870
rect 41921 4868 41977 4870
rect 41681 3834 41737 3836
rect 41761 3834 41817 3836
rect 41841 3834 41897 3836
rect 41921 3834 41977 3836
rect 41681 3782 41707 3834
rect 41707 3782 41737 3834
rect 41761 3782 41771 3834
rect 41771 3782 41817 3834
rect 41841 3782 41887 3834
rect 41887 3782 41897 3834
rect 41921 3782 41951 3834
rect 41951 3782 41977 3834
rect 41681 3780 41737 3782
rect 41761 3780 41817 3782
rect 41841 3780 41897 3782
rect 41921 3780 41977 3782
rect 42062 3440 42118 3496
rect 41326 3304 41382 3360
rect 38750 2896 38806 2952
rect 51862 17434 51918 17436
rect 51942 17434 51998 17436
rect 52022 17434 52078 17436
rect 52102 17434 52158 17436
rect 51862 17382 51888 17434
rect 51888 17382 51918 17434
rect 51942 17382 51952 17434
rect 51952 17382 51998 17434
rect 52022 17382 52068 17434
rect 52068 17382 52078 17434
rect 52102 17382 52132 17434
rect 52132 17382 52158 17434
rect 51862 17380 51918 17382
rect 51942 17380 51998 17382
rect 52022 17380 52078 17382
rect 52102 17380 52158 17382
rect 45190 11620 45246 11656
rect 45190 11600 45192 11620
rect 45192 11600 45244 11620
rect 45244 11600 45246 11620
rect 44178 9016 44234 9072
rect 44178 8200 44234 8256
rect 44454 7248 44510 7304
rect 44362 6740 44364 6760
rect 44364 6740 44416 6760
rect 44416 6740 44418 6760
rect 44362 6704 44418 6740
rect 45374 9016 45430 9072
rect 46294 11872 46350 11928
rect 45742 7828 45744 7848
rect 45744 7828 45796 7848
rect 45796 7828 45798 7848
rect 45742 7792 45798 7828
rect 45190 5752 45246 5808
rect 45650 5772 45706 5808
rect 45650 5752 45652 5772
rect 45652 5752 45704 5772
rect 45704 5752 45706 5772
rect 51862 16346 51918 16348
rect 51942 16346 51998 16348
rect 52022 16346 52078 16348
rect 52102 16346 52158 16348
rect 51862 16294 51888 16346
rect 51888 16294 51918 16346
rect 51942 16294 51952 16346
rect 51952 16294 51998 16346
rect 52022 16294 52068 16346
rect 52068 16294 52078 16346
rect 52102 16294 52132 16346
rect 52132 16294 52158 16346
rect 51862 16292 51918 16294
rect 51942 16292 51998 16294
rect 52022 16292 52078 16294
rect 52102 16292 52158 16294
rect 45926 6432 45982 6488
rect 47306 8744 47362 8800
rect 47306 7384 47362 7440
rect 47306 6840 47362 6896
rect 46754 5480 46810 5536
rect 46754 5072 46810 5128
rect 47490 5208 47546 5264
rect 51862 15258 51918 15260
rect 51942 15258 51998 15260
rect 52022 15258 52078 15260
rect 52102 15258 52158 15260
rect 51862 15206 51888 15258
rect 51888 15206 51918 15258
rect 51942 15206 51952 15258
rect 51952 15206 51998 15258
rect 52022 15206 52068 15258
rect 52068 15206 52078 15258
rect 52102 15206 52132 15258
rect 52132 15206 52158 15258
rect 51862 15204 51918 15206
rect 51942 15204 51998 15206
rect 52022 15204 52078 15206
rect 52102 15204 52158 15206
rect 51862 14170 51918 14172
rect 51942 14170 51998 14172
rect 52022 14170 52078 14172
rect 52102 14170 52158 14172
rect 51862 14118 51888 14170
rect 51888 14118 51918 14170
rect 51942 14118 51952 14170
rect 51952 14118 51998 14170
rect 52022 14118 52068 14170
rect 52068 14118 52078 14170
rect 52102 14118 52132 14170
rect 52132 14118 52158 14170
rect 51862 14116 51918 14118
rect 51942 14116 51998 14118
rect 52022 14116 52078 14118
rect 52102 14116 52158 14118
rect 48686 11620 48742 11656
rect 48686 11600 48688 11620
rect 48688 11600 48740 11620
rect 48740 11600 48742 11620
rect 48134 10512 48190 10568
rect 47950 9036 48006 9072
rect 47950 9016 47952 9036
rect 47952 9016 48004 9036
rect 48004 9016 48006 9036
rect 48502 9016 48558 9072
rect 48410 8744 48466 8800
rect 46938 5072 46994 5128
rect 48318 6840 48374 6896
rect 41681 2746 41737 2748
rect 41761 2746 41817 2748
rect 41841 2746 41897 2748
rect 41921 2746 41977 2748
rect 41681 2694 41707 2746
rect 41707 2694 41737 2746
rect 41761 2694 41771 2746
rect 41771 2694 41817 2746
rect 41841 2694 41887 2746
rect 41887 2694 41897 2746
rect 41921 2694 41951 2746
rect 41951 2694 41977 2746
rect 41681 2692 41737 2694
rect 41761 2692 41817 2694
rect 41841 2692 41897 2694
rect 41921 2692 41977 2694
rect 51862 13082 51918 13084
rect 51942 13082 51998 13084
rect 52022 13082 52078 13084
rect 52102 13082 52158 13084
rect 51862 13030 51888 13082
rect 51888 13030 51918 13082
rect 51942 13030 51952 13082
rect 51952 13030 51998 13082
rect 52022 13030 52068 13082
rect 52068 13030 52078 13082
rect 52102 13030 52132 13082
rect 52132 13030 52158 13082
rect 51862 13028 51918 13030
rect 51942 13028 51998 13030
rect 52022 13028 52078 13030
rect 52102 13028 52158 13030
rect 50250 8608 50306 8664
rect 49330 6740 49332 6760
rect 49332 6740 49384 6760
rect 49384 6740 49386 6760
rect 49330 6704 49386 6740
rect 49514 6196 49516 6216
rect 49516 6196 49568 6216
rect 49568 6196 49570 6216
rect 49514 6160 49570 6196
rect 49330 6024 49386 6080
rect 49422 5908 49478 5944
rect 49422 5888 49424 5908
rect 49424 5888 49476 5908
rect 49476 5888 49478 5908
rect 49238 5752 49294 5808
rect 51862 11994 51918 11996
rect 51942 11994 51998 11996
rect 52022 11994 52078 11996
rect 52102 11994 52158 11996
rect 51862 11942 51888 11994
rect 51888 11942 51918 11994
rect 51942 11942 51952 11994
rect 51952 11942 51998 11994
rect 52022 11942 52068 11994
rect 52068 11942 52078 11994
rect 52102 11942 52132 11994
rect 52132 11942 52158 11994
rect 51862 11940 51918 11942
rect 51942 11940 51998 11942
rect 52022 11940 52078 11942
rect 52102 11940 52158 11942
rect 51262 6860 51318 6896
rect 51262 6840 51264 6860
rect 51264 6840 51316 6860
rect 51316 6840 51318 6860
rect 51262 6432 51318 6488
rect 50710 6296 50766 6352
rect 51170 6316 51226 6352
rect 51170 6296 51172 6316
rect 51172 6296 51224 6316
rect 51224 6296 51226 6316
rect 51862 10906 51918 10908
rect 51942 10906 51998 10908
rect 52022 10906 52078 10908
rect 52102 10906 52158 10908
rect 51862 10854 51888 10906
rect 51888 10854 51918 10906
rect 51942 10854 51952 10906
rect 51952 10854 51998 10906
rect 52022 10854 52068 10906
rect 52068 10854 52078 10906
rect 52102 10854 52132 10906
rect 52132 10854 52158 10906
rect 51862 10852 51918 10854
rect 51942 10852 51998 10854
rect 52022 10852 52078 10854
rect 52102 10852 52158 10854
rect 51862 9818 51918 9820
rect 51942 9818 51998 9820
rect 52022 9818 52078 9820
rect 52102 9818 52158 9820
rect 51862 9766 51888 9818
rect 51888 9766 51918 9818
rect 51942 9766 51952 9818
rect 51952 9766 51998 9818
rect 52022 9766 52068 9818
rect 52068 9766 52078 9818
rect 52102 9766 52132 9818
rect 52132 9766 52158 9818
rect 51862 9764 51918 9766
rect 51942 9764 51998 9766
rect 52022 9764 52078 9766
rect 52102 9764 52158 9766
rect 52918 11600 52974 11656
rect 51862 8730 51918 8732
rect 51942 8730 51998 8732
rect 52022 8730 52078 8732
rect 52102 8730 52158 8732
rect 51862 8678 51888 8730
rect 51888 8678 51918 8730
rect 51942 8678 51952 8730
rect 51952 8678 51998 8730
rect 52022 8678 52068 8730
rect 52068 8678 52078 8730
rect 52102 8678 52132 8730
rect 52132 8678 52158 8730
rect 51862 8676 51918 8678
rect 51942 8676 51998 8678
rect 52022 8676 52078 8678
rect 52102 8676 52158 8678
rect 51862 7642 51918 7644
rect 51942 7642 51998 7644
rect 52022 7642 52078 7644
rect 52102 7642 52158 7644
rect 51862 7590 51888 7642
rect 51888 7590 51918 7642
rect 51942 7590 51952 7642
rect 51952 7590 51998 7642
rect 52022 7590 52068 7642
rect 52068 7590 52078 7642
rect 52102 7590 52132 7642
rect 52132 7590 52158 7642
rect 51862 7588 51918 7590
rect 51942 7588 51998 7590
rect 52022 7588 52078 7590
rect 52102 7588 52158 7590
rect 51862 6554 51918 6556
rect 51942 6554 51998 6556
rect 52022 6554 52078 6556
rect 52102 6554 52158 6556
rect 51862 6502 51888 6554
rect 51888 6502 51918 6554
rect 51942 6502 51952 6554
rect 51952 6502 51998 6554
rect 52022 6502 52068 6554
rect 52068 6502 52078 6554
rect 52102 6502 52132 6554
rect 52132 6502 52158 6554
rect 51862 6500 51918 6502
rect 51942 6500 51998 6502
rect 52022 6500 52078 6502
rect 52102 6500 52158 6502
rect 52274 6160 52330 6216
rect 52182 5752 52238 5808
rect 52458 6704 52514 6760
rect 52918 6604 52920 6624
rect 52920 6604 52972 6624
rect 52972 6604 52974 6624
rect 52918 6568 52974 6604
rect 51862 5466 51918 5468
rect 51942 5466 51998 5468
rect 52022 5466 52078 5468
rect 52102 5466 52158 5468
rect 51862 5414 51888 5466
rect 51888 5414 51918 5466
rect 51942 5414 51952 5466
rect 51952 5414 51998 5466
rect 52022 5414 52068 5466
rect 52068 5414 52078 5466
rect 52102 5414 52132 5466
rect 52132 5414 52158 5466
rect 51862 5412 51918 5414
rect 51942 5412 51998 5414
rect 52022 5412 52078 5414
rect 52102 5412 52158 5414
rect 51862 4378 51918 4380
rect 51942 4378 51998 4380
rect 52022 4378 52078 4380
rect 52102 4378 52158 4380
rect 51862 4326 51888 4378
rect 51888 4326 51918 4378
rect 51942 4326 51952 4378
rect 51952 4326 51998 4378
rect 52022 4326 52068 4378
rect 52068 4326 52078 4378
rect 52102 4326 52132 4378
rect 52132 4326 52158 4378
rect 51862 4324 51918 4326
rect 51942 4324 51998 4326
rect 52022 4324 52078 4326
rect 52102 4324 52158 4326
rect 53654 8372 53656 8392
rect 53656 8372 53708 8392
rect 53708 8372 53710 8392
rect 53654 8336 53710 8372
rect 53746 6568 53802 6624
rect 53746 6296 53802 6352
rect 53562 5888 53618 5944
rect 54022 6840 54078 6896
rect 53930 6316 53986 6352
rect 53930 6296 53932 6316
rect 53932 6296 53984 6316
rect 53984 6296 53986 6316
rect 54666 6024 54722 6080
rect 53102 3576 53158 3632
rect 48686 3168 48742 3224
rect 51862 3290 51918 3292
rect 51942 3290 51998 3292
rect 52022 3290 52078 3292
rect 52102 3290 52158 3292
rect 51862 3238 51888 3290
rect 51888 3238 51918 3290
rect 51942 3238 51952 3290
rect 51952 3238 51998 3290
rect 52022 3238 52068 3290
rect 52068 3238 52078 3290
rect 52102 3238 52132 3290
rect 52132 3238 52158 3290
rect 51862 3236 51918 3238
rect 51942 3236 51998 3238
rect 52022 3236 52078 3238
rect 52102 3236 52158 3238
rect 52458 2896 52514 2952
rect 51862 2202 51918 2204
rect 51942 2202 51998 2204
rect 52022 2202 52078 2204
rect 52102 2202 52158 2204
rect 51862 2150 51888 2202
rect 51888 2150 51918 2202
rect 51942 2150 51952 2202
rect 51952 2150 51998 2202
rect 52022 2150 52068 2202
rect 52068 2150 52078 2202
rect 52102 2150 52132 2202
rect 52132 2150 52158 2202
rect 51862 2148 51918 2150
rect 51942 2148 51998 2150
rect 52022 2148 52078 2150
rect 52102 2148 52158 2150
rect 54022 3576 54078 3632
rect 55862 8472 55918 8528
rect 55126 6296 55182 6352
rect 57058 9036 57114 9072
rect 57058 9016 57060 9036
rect 57060 9016 57112 9036
rect 57112 9016 57114 9036
rect 56690 8880 56746 8936
rect 57242 7928 57298 7984
rect 58714 8880 58770 8936
rect 56506 3984 56562 4040
rect 55586 3032 55642 3088
rect 55586 2932 55588 2952
rect 55588 2932 55640 2952
rect 55640 2932 55642 2952
rect 55586 2896 55642 2932
rect 56874 3596 56930 3632
rect 56874 3576 56876 3596
rect 56876 3576 56928 3596
rect 56928 3576 56930 3596
<< metal3 >>
rect 0 18594 800 18624
rect 3325 18594 3391 18597
rect 0 18592 3391 18594
rect 0 18536 3330 18592
rect 3386 18536 3391 18592
rect 0 18534 3391 18536
rect 0 18504 800 18534
rect 3325 18531 3391 18534
rect 11125 17440 11445 17441
rect 11125 17376 11133 17440
rect 11197 17376 11213 17440
rect 11277 17376 11293 17440
rect 11357 17376 11373 17440
rect 11437 17376 11445 17440
rect 11125 17375 11445 17376
rect 31488 17440 31808 17441
rect 31488 17376 31496 17440
rect 31560 17376 31576 17440
rect 31640 17376 31656 17440
rect 31720 17376 31736 17440
rect 31800 17376 31808 17440
rect 31488 17375 31808 17376
rect 51850 17440 52170 17441
rect 51850 17376 51858 17440
rect 51922 17376 51938 17440
rect 52002 17376 52018 17440
rect 52082 17376 52098 17440
rect 52162 17376 52170 17440
rect 51850 17375 52170 17376
rect 21306 16896 21626 16897
rect 21306 16832 21314 16896
rect 21378 16832 21394 16896
rect 21458 16832 21474 16896
rect 21538 16832 21554 16896
rect 21618 16832 21626 16896
rect 21306 16831 21626 16832
rect 41669 16896 41989 16897
rect 41669 16832 41677 16896
rect 41741 16832 41757 16896
rect 41821 16832 41837 16896
rect 41901 16832 41917 16896
rect 41981 16832 41989 16896
rect 41669 16831 41989 16832
rect 0 16418 800 16448
rect 3049 16418 3115 16421
rect 0 16416 3115 16418
rect 0 16360 3054 16416
rect 3110 16360 3115 16416
rect 0 16358 3115 16360
rect 0 16328 800 16358
rect 3049 16355 3115 16358
rect 11125 16352 11445 16353
rect 11125 16288 11133 16352
rect 11197 16288 11213 16352
rect 11277 16288 11293 16352
rect 11357 16288 11373 16352
rect 11437 16288 11445 16352
rect 11125 16287 11445 16288
rect 31488 16352 31808 16353
rect 31488 16288 31496 16352
rect 31560 16288 31576 16352
rect 31640 16288 31656 16352
rect 31720 16288 31736 16352
rect 31800 16288 31808 16352
rect 31488 16287 31808 16288
rect 51850 16352 52170 16353
rect 51850 16288 51858 16352
rect 51922 16288 51938 16352
rect 52002 16288 52018 16352
rect 52082 16288 52098 16352
rect 52162 16288 52170 16352
rect 51850 16287 52170 16288
rect 21306 15808 21626 15809
rect 21306 15744 21314 15808
rect 21378 15744 21394 15808
rect 21458 15744 21474 15808
rect 21538 15744 21554 15808
rect 21618 15744 21626 15808
rect 21306 15743 21626 15744
rect 41669 15808 41989 15809
rect 41669 15744 41677 15808
rect 41741 15744 41757 15808
rect 41821 15744 41837 15808
rect 41901 15744 41917 15808
rect 41981 15744 41989 15808
rect 41669 15743 41989 15744
rect 11125 15264 11445 15265
rect 11125 15200 11133 15264
rect 11197 15200 11213 15264
rect 11277 15200 11293 15264
rect 11357 15200 11373 15264
rect 11437 15200 11445 15264
rect 11125 15199 11445 15200
rect 31488 15264 31808 15265
rect 31488 15200 31496 15264
rect 31560 15200 31576 15264
rect 31640 15200 31656 15264
rect 31720 15200 31736 15264
rect 31800 15200 31808 15264
rect 31488 15199 31808 15200
rect 51850 15264 52170 15265
rect 51850 15200 51858 15264
rect 51922 15200 51938 15264
rect 52002 15200 52018 15264
rect 52082 15200 52098 15264
rect 52162 15200 52170 15264
rect 51850 15199 52170 15200
rect 21306 14720 21626 14721
rect 21306 14656 21314 14720
rect 21378 14656 21394 14720
rect 21458 14656 21474 14720
rect 21538 14656 21554 14720
rect 21618 14656 21626 14720
rect 21306 14655 21626 14656
rect 41669 14720 41989 14721
rect 41669 14656 41677 14720
rect 41741 14656 41757 14720
rect 41821 14656 41837 14720
rect 41901 14656 41917 14720
rect 41981 14656 41989 14720
rect 41669 14655 41989 14656
rect 0 14242 800 14272
rect 4061 14242 4127 14245
rect 0 14240 4127 14242
rect 0 14184 4066 14240
rect 4122 14184 4127 14240
rect 0 14182 4127 14184
rect 0 14152 800 14182
rect 4061 14179 4127 14182
rect 11125 14176 11445 14177
rect 11125 14112 11133 14176
rect 11197 14112 11213 14176
rect 11277 14112 11293 14176
rect 11357 14112 11373 14176
rect 11437 14112 11445 14176
rect 11125 14111 11445 14112
rect 31488 14176 31808 14177
rect 31488 14112 31496 14176
rect 31560 14112 31576 14176
rect 31640 14112 31656 14176
rect 31720 14112 31736 14176
rect 31800 14112 31808 14176
rect 31488 14111 31808 14112
rect 51850 14176 52170 14177
rect 51850 14112 51858 14176
rect 51922 14112 51938 14176
rect 52002 14112 52018 14176
rect 52082 14112 52098 14176
rect 52162 14112 52170 14176
rect 51850 14111 52170 14112
rect 21306 13632 21626 13633
rect 21306 13568 21314 13632
rect 21378 13568 21394 13632
rect 21458 13568 21474 13632
rect 21538 13568 21554 13632
rect 21618 13568 21626 13632
rect 21306 13567 21626 13568
rect 41669 13632 41989 13633
rect 41669 13568 41677 13632
rect 41741 13568 41757 13632
rect 41821 13568 41837 13632
rect 41901 13568 41917 13632
rect 41981 13568 41989 13632
rect 41669 13567 41989 13568
rect 10961 13562 11027 13565
rect 16573 13562 16639 13565
rect 10961 13560 16639 13562
rect 10961 13504 10966 13560
rect 11022 13504 16578 13560
rect 16634 13504 16639 13560
rect 10961 13502 16639 13504
rect 10961 13499 11027 13502
rect 16573 13499 16639 13502
rect 19425 13426 19491 13429
rect 23013 13426 23079 13429
rect 19425 13424 23079 13426
rect 19425 13368 19430 13424
rect 19486 13368 23018 13424
rect 23074 13368 23079 13424
rect 19425 13366 23079 13368
rect 19425 13363 19491 13366
rect 23013 13363 23079 13366
rect 10777 13290 10843 13293
rect 15285 13290 15351 13293
rect 19057 13290 19123 13293
rect 10777 13288 19123 13290
rect 10777 13232 10782 13288
rect 10838 13232 15290 13288
rect 15346 13232 19062 13288
rect 19118 13232 19123 13288
rect 10777 13230 19123 13232
rect 10777 13227 10843 13230
rect 15285 13227 15351 13230
rect 19057 13227 19123 13230
rect 20345 13154 20411 13157
rect 27061 13154 27127 13157
rect 20345 13152 27127 13154
rect 20345 13096 20350 13152
rect 20406 13096 27066 13152
rect 27122 13096 27127 13152
rect 20345 13094 27127 13096
rect 20345 13091 20411 13094
rect 27061 13091 27127 13094
rect 11125 13088 11445 13089
rect 11125 13024 11133 13088
rect 11197 13024 11213 13088
rect 11277 13024 11293 13088
rect 11357 13024 11373 13088
rect 11437 13024 11445 13088
rect 11125 13023 11445 13024
rect 31488 13088 31808 13089
rect 31488 13024 31496 13088
rect 31560 13024 31576 13088
rect 31640 13024 31656 13088
rect 31720 13024 31736 13088
rect 31800 13024 31808 13088
rect 31488 13023 31808 13024
rect 51850 13088 52170 13089
rect 51850 13024 51858 13088
rect 51922 13024 51938 13088
rect 52002 13024 52018 13088
rect 52082 13024 52098 13088
rect 52162 13024 52170 13088
rect 51850 13023 52170 13024
rect 20437 13018 20503 13021
rect 26877 13018 26943 13021
rect 20437 13016 26943 13018
rect 20437 12960 20442 13016
rect 20498 12960 26882 13016
rect 26938 12960 26943 13016
rect 20437 12958 26943 12960
rect 20437 12955 20503 12958
rect 26877 12955 26943 12958
rect 22645 12882 22711 12885
rect 27705 12882 27771 12885
rect 22645 12880 27771 12882
rect 22645 12824 22650 12880
rect 22706 12824 27710 12880
rect 27766 12824 27771 12880
rect 22645 12822 27771 12824
rect 22645 12819 22711 12822
rect 27705 12819 27771 12822
rect 33869 12882 33935 12885
rect 36077 12882 36143 12885
rect 33869 12880 36143 12882
rect 33869 12824 33874 12880
rect 33930 12824 36082 12880
rect 36138 12824 36143 12880
rect 33869 12822 36143 12824
rect 33869 12819 33935 12822
rect 36077 12819 36143 12822
rect 29361 12746 29427 12749
rect 34237 12746 34303 12749
rect 29361 12744 34303 12746
rect 29361 12688 29366 12744
rect 29422 12688 34242 12744
rect 34298 12688 34303 12744
rect 29361 12686 34303 12688
rect 29361 12683 29427 12686
rect 34237 12683 34303 12686
rect 26325 12610 26391 12613
rect 27889 12610 27955 12613
rect 26325 12608 27955 12610
rect 26325 12552 26330 12608
rect 26386 12552 27894 12608
rect 27950 12552 27955 12608
rect 26325 12550 27955 12552
rect 26325 12547 26391 12550
rect 27889 12547 27955 12550
rect 21306 12544 21626 12545
rect 21306 12480 21314 12544
rect 21378 12480 21394 12544
rect 21458 12480 21474 12544
rect 21538 12480 21554 12544
rect 21618 12480 21626 12544
rect 21306 12479 21626 12480
rect 41669 12544 41989 12545
rect 41669 12480 41677 12544
rect 41741 12480 41757 12544
rect 41821 12480 41837 12544
rect 41901 12480 41917 12544
rect 41981 12480 41989 12544
rect 41669 12479 41989 12480
rect 30005 12474 30071 12477
rect 37365 12474 37431 12477
rect 30005 12472 37431 12474
rect 30005 12416 30010 12472
rect 30066 12416 37370 12472
rect 37426 12416 37431 12472
rect 30005 12414 37431 12416
rect 30005 12411 30071 12414
rect 37365 12411 37431 12414
rect 9857 12338 9923 12341
rect 17769 12338 17835 12341
rect 9857 12336 17835 12338
rect 9857 12280 9862 12336
rect 9918 12280 17774 12336
rect 17830 12280 17835 12336
rect 9857 12278 17835 12280
rect 9857 12275 9923 12278
rect 17769 12275 17835 12278
rect 30465 12202 30531 12205
rect 31201 12202 31267 12205
rect 30465 12200 31267 12202
rect 30465 12144 30470 12200
rect 30526 12144 31206 12200
rect 31262 12144 31267 12200
rect 30465 12142 31267 12144
rect 30465 12139 30531 12142
rect 31201 12139 31267 12142
rect 0 12066 800 12096
rect 3509 12066 3575 12069
rect 0 12064 3575 12066
rect 0 12008 3514 12064
rect 3570 12008 3575 12064
rect 0 12006 3575 12008
rect 0 11976 800 12006
rect 3509 12003 3575 12006
rect 11125 12000 11445 12001
rect 11125 11936 11133 12000
rect 11197 11936 11213 12000
rect 11277 11936 11293 12000
rect 11357 11936 11373 12000
rect 11437 11936 11445 12000
rect 11125 11935 11445 11936
rect 31488 12000 31808 12001
rect 31488 11936 31496 12000
rect 31560 11936 31576 12000
rect 31640 11936 31656 12000
rect 31720 11936 31736 12000
rect 31800 11936 31808 12000
rect 31488 11935 31808 11936
rect 51850 12000 52170 12001
rect 51850 11936 51858 12000
rect 51922 11936 51938 12000
rect 52002 11936 52018 12000
rect 52082 11936 52098 12000
rect 52162 11936 52170 12000
rect 51850 11935 52170 11936
rect 12893 11930 12959 11933
rect 16389 11930 16455 11933
rect 18873 11930 18939 11933
rect 12893 11928 18939 11930
rect 12893 11872 12898 11928
rect 12954 11872 16394 11928
rect 16450 11872 18878 11928
rect 18934 11872 18939 11928
rect 12893 11870 18939 11872
rect 12893 11867 12959 11870
rect 16389 11867 16455 11870
rect 18873 11867 18939 11870
rect 39665 11930 39731 11933
rect 46289 11930 46355 11933
rect 39665 11928 46355 11930
rect 39665 11872 39670 11928
rect 39726 11872 46294 11928
rect 46350 11872 46355 11928
rect 39665 11870 46355 11872
rect 39665 11867 39731 11870
rect 46289 11867 46355 11870
rect 12341 11794 12407 11797
rect 13261 11794 13327 11797
rect 12341 11792 13327 11794
rect 12341 11736 12346 11792
rect 12402 11736 13266 11792
rect 13322 11736 13327 11792
rect 12341 11734 13327 11736
rect 12341 11731 12407 11734
rect 13261 11731 13327 11734
rect 20805 11794 20871 11797
rect 23749 11794 23815 11797
rect 20805 11792 23815 11794
rect 20805 11736 20810 11792
rect 20866 11736 23754 11792
rect 23810 11736 23815 11792
rect 20805 11734 23815 11736
rect 20805 11731 20871 11734
rect 23749 11731 23815 11734
rect 11237 11658 11303 11661
rect 13353 11658 13419 11661
rect 11237 11656 13419 11658
rect 11237 11600 11242 11656
rect 11298 11600 13358 11656
rect 13414 11600 13419 11656
rect 11237 11598 13419 11600
rect 11237 11595 11303 11598
rect 13353 11595 13419 11598
rect 41229 11658 41295 11661
rect 45185 11658 45251 11661
rect 41229 11656 45251 11658
rect 41229 11600 41234 11656
rect 41290 11600 45190 11656
rect 45246 11600 45251 11656
rect 41229 11598 45251 11600
rect 41229 11595 41295 11598
rect 45185 11595 45251 11598
rect 48681 11658 48747 11661
rect 52913 11658 52979 11661
rect 48681 11656 52979 11658
rect 48681 11600 48686 11656
rect 48742 11600 52918 11656
rect 52974 11600 52979 11656
rect 48681 11598 52979 11600
rect 48681 11595 48747 11598
rect 52913 11595 52979 11598
rect 13169 11522 13235 11525
rect 18781 11522 18847 11525
rect 13169 11520 18847 11522
rect 13169 11464 13174 11520
rect 13230 11464 18786 11520
rect 18842 11464 18847 11520
rect 13169 11462 18847 11464
rect 13169 11459 13235 11462
rect 18781 11459 18847 11462
rect 21306 11456 21626 11457
rect 21306 11392 21314 11456
rect 21378 11392 21394 11456
rect 21458 11392 21474 11456
rect 21538 11392 21554 11456
rect 21618 11392 21626 11456
rect 21306 11391 21626 11392
rect 41669 11456 41989 11457
rect 41669 11392 41677 11456
rect 41741 11392 41757 11456
rect 41821 11392 41837 11456
rect 41901 11392 41917 11456
rect 41981 11392 41989 11456
rect 41669 11391 41989 11392
rect 10777 11250 10843 11253
rect 14549 11250 14615 11253
rect 10777 11248 14615 11250
rect 10777 11192 10782 11248
rect 10838 11192 14554 11248
rect 14610 11192 14615 11248
rect 10777 11190 14615 11192
rect 10777 11187 10843 11190
rect 14549 11187 14615 11190
rect 21081 11250 21147 11253
rect 27797 11250 27863 11253
rect 21081 11248 27863 11250
rect 21081 11192 21086 11248
rect 21142 11192 27802 11248
rect 27858 11192 27863 11248
rect 21081 11190 27863 11192
rect 21081 11187 21147 11190
rect 27797 11187 27863 11190
rect 20897 11114 20963 11117
rect 24945 11114 25011 11117
rect 20897 11112 25011 11114
rect 20897 11056 20902 11112
rect 20958 11056 24950 11112
rect 25006 11056 25011 11112
rect 20897 11054 25011 11056
rect 20897 11051 20963 11054
rect 24945 11051 25011 11054
rect 11125 10912 11445 10913
rect 11125 10848 11133 10912
rect 11197 10848 11213 10912
rect 11277 10848 11293 10912
rect 11357 10848 11373 10912
rect 11437 10848 11445 10912
rect 11125 10847 11445 10848
rect 31488 10912 31808 10913
rect 31488 10848 31496 10912
rect 31560 10848 31576 10912
rect 31640 10848 31656 10912
rect 31720 10848 31736 10912
rect 31800 10848 31808 10912
rect 31488 10847 31808 10848
rect 51850 10912 52170 10913
rect 51850 10848 51858 10912
rect 51922 10848 51938 10912
rect 52002 10848 52018 10912
rect 52082 10848 52098 10912
rect 52162 10848 52170 10912
rect 51850 10847 52170 10848
rect 11605 10842 11671 10845
rect 20897 10842 20963 10845
rect 11605 10840 20963 10842
rect 11605 10784 11610 10840
rect 11666 10784 20902 10840
rect 20958 10784 20963 10840
rect 11605 10782 20963 10784
rect 11605 10779 11671 10782
rect 20897 10779 20963 10782
rect 8753 10570 8819 10573
rect 9213 10570 9279 10573
rect 28625 10570 28691 10573
rect 48129 10570 48195 10573
rect 8753 10568 48195 10570
rect 8753 10512 8758 10568
rect 8814 10512 9218 10568
rect 9274 10512 28630 10568
rect 28686 10512 48134 10568
rect 48190 10512 48195 10568
rect 8753 10510 48195 10512
rect 8753 10507 8819 10510
rect 9213 10507 9279 10510
rect 28625 10507 28691 10510
rect 48129 10507 48195 10510
rect 21306 10368 21626 10369
rect 21306 10304 21314 10368
rect 21378 10304 21394 10368
rect 21458 10304 21474 10368
rect 21538 10304 21554 10368
rect 21618 10304 21626 10368
rect 21306 10303 21626 10304
rect 41669 10368 41989 10369
rect 41669 10304 41677 10368
rect 41741 10304 41757 10368
rect 41821 10304 41837 10368
rect 41901 10304 41917 10368
rect 41981 10304 41989 10368
rect 41669 10303 41989 10304
rect 19333 10026 19399 10029
rect 20989 10026 21055 10029
rect 19333 10024 21055 10026
rect 19333 9968 19338 10024
rect 19394 9968 20994 10024
rect 21050 9968 21055 10024
rect 19333 9966 21055 9968
rect 19333 9963 19399 9966
rect 20989 9963 21055 9966
rect 0 9890 800 9920
rect 2773 9890 2839 9893
rect 0 9888 2839 9890
rect 0 9832 2778 9888
rect 2834 9832 2839 9888
rect 0 9830 2839 9832
rect 0 9800 800 9830
rect 2773 9827 2839 9830
rect 11125 9824 11445 9825
rect 11125 9760 11133 9824
rect 11197 9760 11213 9824
rect 11277 9760 11293 9824
rect 11357 9760 11373 9824
rect 11437 9760 11445 9824
rect 11125 9759 11445 9760
rect 31488 9824 31808 9825
rect 31488 9760 31496 9824
rect 31560 9760 31576 9824
rect 31640 9760 31656 9824
rect 31720 9760 31736 9824
rect 31800 9760 31808 9824
rect 31488 9759 31808 9760
rect 51850 9824 52170 9825
rect 51850 9760 51858 9824
rect 51922 9760 51938 9824
rect 52002 9760 52018 9824
rect 52082 9760 52098 9824
rect 52162 9760 52170 9824
rect 51850 9759 52170 9760
rect 20805 9754 20871 9757
rect 31293 9754 31359 9757
rect 20805 9752 31359 9754
rect 20805 9696 20810 9752
rect 20866 9696 31298 9752
rect 31354 9696 31359 9752
rect 20805 9694 31359 9696
rect 20805 9691 20871 9694
rect 31293 9691 31359 9694
rect 19609 9618 19675 9621
rect 23749 9618 23815 9621
rect 25221 9618 25287 9621
rect 19609 9616 25287 9618
rect 19609 9560 19614 9616
rect 19670 9560 23754 9616
rect 23810 9560 25226 9616
rect 25282 9560 25287 9616
rect 19609 9558 25287 9560
rect 19609 9555 19675 9558
rect 23749 9555 23815 9558
rect 25221 9555 25287 9558
rect 37273 9618 37339 9621
rect 41413 9618 41479 9621
rect 37273 9616 41479 9618
rect 37273 9560 37278 9616
rect 37334 9560 41418 9616
rect 41474 9560 41479 9616
rect 37273 9558 41479 9560
rect 37273 9555 37339 9558
rect 41413 9555 41479 9558
rect 21306 9280 21626 9281
rect 21306 9216 21314 9280
rect 21378 9216 21394 9280
rect 21458 9216 21474 9280
rect 21538 9216 21554 9280
rect 21618 9216 21626 9280
rect 21306 9215 21626 9216
rect 41669 9280 41989 9281
rect 41669 9216 41677 9280
rect 41741 9216 41757 9280
rect 41821 9216 41837 9280
rect 41901 9216 41917 9280
rect 41981 9216 41989 9280
rect 41669 9215 41989 9216
rect 12341 9074 12407 9077
rect 17953 9074 18019 9077
rect 12341 9072 18019 9074
rect 12341 9016 12346 9072
rect 12402 9016 17958 9072
rect 18014 9016 18019 9072
rect 12341 9014 18019 9016
rect 12341 9011 12407 9014
rect 17953 9011 18019 9014
rect 20253 9074 20319 9077
rect 21541 9074 21607 9077
rect 27705 9074 27771 9077
rect 20253 9072 27771 9074
rect 20253 9016 20258 9072
rect 20314 9016 21546 9072
rect 21602 9016 27710 9072
rect 27766 9016 27771 9072
rect 20253 9014 27771 9016
rect 20253 9011 20319 9014
rect 21541 9011 21607 9014
rect 27705 9011 27771 9014
rect 44173 9074 44239 9077
rect 45369 9074 45435 9077
rect 47945 9074 48011 9077
rect 44173 9072 48011 9074
rect 44173 9016 44178 9072
rect 44234 9016 45374 9072
rect 45430 9016 47950 9072
rect 48006 9016 48011 9072
rect 44173 9014 48011 9016
rect 44173 9011 44239 9014
rect 45369 9011 45435 9014
rect 47945 9011 48011 9014
rect 48497 9074 48563 9077
rect 57053 9074 57119 9077
rect 48497 9072 57119 9074
rect 48497 9016 48502 9072
rect 48558 9016 57058 9072
rect 57114 9016 57119 9072
rect 48497 9014 57119 9016
rect 48497 9011 48563 9014
rect 57053 9011 57119 9014
rect 17769 8938 17835 8941
rect 20897 8938 20963 8941
rect 17769 8936 20963 8938
rect 17769 8880 17774 8936
rect 17830 8880 20902 8936
rect 20958 8880 20963 8936
rect 17769 8878 20963 8880
rect 17769 8875 17835 8878
rect 20897 8875 20963 8878
rect 56685 8938 56751 8941
rect 58709 8938 58775 8941
rect 56685 8936 58775 8938
rect 56685 8880 56690 8936
rect 56746 8880 58714 8936
rect 58770 8880 58775 8936
rect 56685 8878 58775 8880
rect 56685 8875 56751 8878
rect 58709 8875 58775 8878
rect 47301 8802 47367 8805
rect 48405 8802 48471 8805
rect 47301 8800 48471 8802
rect 47301 8744 47306 8800
rect 47362 8744 48410 8800
rect 48466 8744 48471 8800
rect 47301 8742 48471 8744
rect 47301 8739 47367 8742
rect 48405 8739 48471 8742
rect 11125 8736 11445 8737
rect 11125 8672 11133 8736
rect 11197 8672 11213 8736
rect 11277 8672 11293 8736
rect 11357 8672 11373 8736
rect 11437 8672 11445 8736
rect 11125 8671 11445 8672
rect 31488 8736 31808 8737
rect 31488 8672 31496 8736
rect 31560 8672 31576 8736
rect 31640 8672 31656 8736
rect 31720 8672 31736 8736
rect 31800 8672 31808 8736
rect 31488 8671 31808 8672
rect 51850 8736 52170 8737
rect 51850 8672 51858 8736
rect 51922 8672 51938 8736
rect 52002 8672 52018 8736
rect 52082 8672 52098 8736
rect 52162 8672 52170 8736
rect 51850 8671 52170 8672
rect 20713 8666 20779 8669
rect 22553 8666 22619 8669
rect 20713 8664 22619 8666
rect 20713 8608 20718 8664
rect 20774 8608 22558 8664
rect 22614 8608 22619 8664
rect 20713 8606 22619 8608
rect 20713 8603 20779 8606
rect 22553 8603 22619 8606
rect 42149 8666 42215 8669
rect 50245 8666 50311 8669
rect 42149 8664 50311 8666
rect 42149 8608 42154 8664
rect 42210 8608 50250 8664
rect 50306 8608 50311 8664
rect 42149 8606 50311 8608
rect 42149 8603 42215 8606
rect 50245 8603 50311 8606
rect 20161 8530 20227 8533
rect 22001 8530 22067 8533
rect 20161 8528 22067 8530
rect 20161 8472 20166 8528
rect 20222 8472 22006 8528
rect 22062 8472 22067 8528
rect 20161 8470 22067 8472
rect 20161 8467 20227 8470
rect 22001 8467 22067 8470
rect 31845 8530 31911 8533
rect 32121 8530 32187 8533
rect 55857 8530 55923 8533
rect 31845 8528 55923 8530
rect 31845 8472 31850 8528
rect 31906 8472 32126 8528
rect 32182 8472 55862 8528
rect 55918 8472 55923 8528
rect 31845 8470 55923 8472
rect 31845 8467 31911 8470
rect 32121 8467 32187 8470
rect 55857 8467 55923 8470
rect 21817 8394 21883 8397
rect 27153 8394 27219 8397
rect 21817 8392 27219 8394
rect 21817 8336 21822 8392
rect 21878 8336 27158 8392
rect 27214 8336 27219 8392
rect 21817 8334 27219 8336
rect 21817 8331 21883 8334
rect 27153 8331 27219 8334
rect 40953 8394 41019 8397
rect 41229 8394 41295 8397
rect 53649 8394 53715 8397
rect 40953 8392 53715 8394
rect 40953 8336 40958 8392
rect 41014 8336 41234 8392
rect 41290 8336 53654 8392
rect 53710 8336 53715 8392
rect 40953 8334 53715 8336
rect 40953 8331 41019 8334
rect 41229 8331 41295 8334
rect 53649 8331 53715 8334
rect 42149 8258 42215 8261
rect 44173 8258 44239 8261
rect 42149 8256 44239 8258
rect 42149 8200 42154 8256
rect 42210 8200 44178 8256
rect 44234 8200 44239 8256
rect 42149 8198 44239 8200
rect 42149 8195 42215 8198
rect 44173 8195 44239 8198
rect 21306 8192 21626 8193
rect 21306 8128 21314 8192
rect 21378 8128 21394 8192
rect 21458 8128 21474 8192
rect 21538 8128 21554 8192
rect 21618 8128 21626 8192
rect 21306 8127 21626 8128
rect 41669 8192 41989 8193
rect 41669 8128 41677 8192
rect 41741 8128 41757 8192
rect 41821 8128 41837 8192
rect 41901 8128 41917 8192
rect 41981 8128 41989 8192
rect 41669 8127 41989 8128
rect 12617 7986 12683 7989
rect 17861 7986 17927 7989
rect 12617 7984 17927 7986
rect 12617 7928 12622 7984
rect 12678 7928 17866 7984
rect 17922 7928 17927 7984
rect 12617 7926 17927 7928
rect 12617 7923 12683 7926
rect 17861 7923 17927 7926
rect 32213 7986 32279 7989
rect 32949 7986 33015 7989
rect 57237 7986 57303 7989
rect 32213 7984 57303 7986
rect 32213 7928 32218 7984
rect 32274 7928 32954 7984
rect 33010 7928 57242 7984
rect 57298 7928 57303 7984
rect 32213 7926 57303 7928
rect 32213 7923 32279 7926
rect 32949 7923 33015 7926
rect 57237 7923 57303 7926
rect 20437 7850 20503 7853
rect 22645 7850 22711 7853
rect 45737 7850 45803 7853
rect 20437 7848 45803 7850
rect 20437 7792 20442 7848
rect 20498 7792 22650 7848
rect 22706 7792 45742 7848
rect 45798 7792 45803 7848
rect 20437 7790 45803 7792
rect 20437 7787 20503 7790
rect 22645 7787 22711 7790
rect 45737 7787 45803 7790
rect 0 7714 800 7744
rect 3049 7714 3115 7717
rect 0 7712 3115 7714
rect 0 7656 3054 7712
rect 3110 7656 3115 7712
rect 0 7654 3115 7656
rect 0 7624 800 7654
rect 3049 7651 3115 7654
rect 11125 7648 11445 7649
rect 11125 7584 11133 7648
rect 11197 7584 11213 7648
rect 11277 7584 11293 7648
rect 11357 7584 11373 7648
rect 11437 7584 11445 7648
rect 11125 7583 11445 7584
rect 31488 7648 31808 7649
rect 31488 7584 31496 7648
rect 31560 7584 31576 7648
rect 31640 7584 31656 7648
rect 31720 7584 31736 7648
rect 31800 7584 31808 7648
rect 31488 7583 31808 7584
rect 51850 7648 52170 7649
rect 51850 7584 51858 7648
rect 51922 7584 51938 7648
rect 52002 7584 52018 7648
rect 52082 7584 52098 7648
rect 52162 7584 52170 7648
rect 51850 7583 52170 7584
rect 40861 7442 40927 7445
rect 47301 7442 47367 7445
rect 40861 7440 47367 7442
rect 40861 7384 40866 7440
rect 40922 7384 47306 7440
rect 47362 7384 47367 7440
rect 40861 7382 47367 7384
rect 40861 7379 40927 7382
rect 47301 7379 47367 7382
rect 32857 7306 32923 7309
rect 44449 7306 44515 7309
rect 32857 7304 44515 7306
rect 32857 7248 32862 7304
rect 32918 7248 44454 7304
rect 44510 7248 44515 7304
rect 32857 7246 44515 7248
rect 32857 7243 32923 7246
rect 44449 7243 44515 7246
rect 30189 7170 30255 7173
rect 35985 7170 36051 7173
rect 30189 7168 36051 7170
rect 30189 7112 30194 7168
rect 30250 7112 35990 7168
rect 36046 7112 36051 7168
rect 30189 7110 36051 7112
rect 30189 7107 30255 7110
rect 35985 7107 36051 7110
rect 38561 7170 38627 7173
rect 38745 7170 38811 7173
rect 38561 7168 38811 7170
rect 38561 7112 38566 7168
rect 38622 7112 38750 7168
rect 38806 7112 38811 7168
rect 38561 7110 38811 7112
rect 38561 7107 38627 7110
rect 38745 7107 38811 7110
rect 21306 7104 21626 7105
rect 21306 7040 21314 7104
rect 21378 7040 21394 7104
rect 21458 7040 21474 7104
rect 21538 7040 21554 7104
rect 21618 7040 21626 7104
rect 21306 7039 21626 7040
rect 41669 7104 41989 7105
rect 41669 7040 41677 7104
rect 41741 7040 41757 7104
rect 41821 7040 41837 7104
rect 41901 7040 41917 7104
rect 41981 7040 41989 7104
rect 41669 7039 41989 7040
rect 28073 7034 28139 7037
rect 32029 7034 32095 7037
rect 28073 7032 32095 7034
rect 28073 6976 28078 7032
rect 28134 6976 32034 7032
rect 32090 6976 32095 7032
rect 28073 6974 32095 6976
rect 28073 6971 28139 6974
rect 32029 6971 32095 6974
rect 35709 7034 35775 7037
rect 41229 7034 41295 7037
rect 35709 7032 41295 7034
rect 35709 6976 35714 7032
rect 35770 6976 41234 7032
rect 41290 6976 41295 7032
rect 35709 6974 41295 6976
rect 35709 6971 35775 6974
rect 41229 6971 41295 6974
rect 1853 6898 1919 6901
rect 47301 6898 47367 6901
rect 1853 6896 47367 6898
rect 1853 6840 1858 6896
rect 1914 6840 47306 6896
rect 47362 6840 47367 6896
rect 1853 6838 47367 6840
rect 1853 6835 1919 6838
rect 47301 6835 47367 6838
rect 48313 6898 48379 6901
rect 51257 6898 51323 6901
rect 54017 6898 54083 6901
rect 48313 6896 54083 6898
rect 48313 6840 48318 6896
rect 48374 6840 51262 6896
rect 51318 6840 54022 6896
rect 54078 6840 54083 6896
rect 48313 6838 54083 6840
rect 48313 6835 48379 6838
rect 51257 6835 51323 6838
rect 54017 6835 54083 6838
rect 20989 6762 21055 6765
rect 32765 6762 32831 6765
rect 20989 6760 32831 6762
rect 20989 6704 20994 6760
rect 21050 6704 32770 6760
rect 32826 6704 32831 6760
rect 20989 6702 32831 6704
rect 20989 6699 21055 6702
rect 32765 6699 32831 6702
rect 37273 6762 37339 6765
rect 44357 6762 44423 6765
rect 37273 6760 44423 6762
rect 37273 6704 37278 6760
rect 37334 6704 44362 6760
rect 44418 6704 44423 6760
rect 37273 6702 44423 6704
rect 37273 6699 37339 6702
rect 44357 6699 44423 6702
rect 49325 6762 49391 6765
rect 52453 6762 52519 6765
rect 49325 6760 52519 6762
rect 49325 6704 49330 6760
rect 49386 6704 52458 6760
rect 52514 6704 52519 6760
rect 49325 6702 52519 6704
rect 49325 6699 49391 6702
rect 52453 6699 52519 6702
rect 52913 6626 52979 6629
rect 53741 6626 53807 6629
rect 52913 6624 53807 6626
rect 52913 6568 52918 6624
rect 52974 6568 53746 6624
rect 53802 6568 53807 6624
rect 52913 6566 53807 6568
rect 52913 6563 52979 6566
rect 53741 6563 53807 6566
rect 11125 6560 11445 6561
rect 11125 6496 11133 6560
rect 11197 6496 11213 6560
rect 11277 6496 11293 6560
rect 11357 6496 11373 6560
rect 11437 6496 11445 6560
rect 11125 6495 11445 6496
rect 31488 6560 31808 6561
rect 31488 6496 31496 6560
rect 31560 6496 31576 6560
rect 31640 6496 31656 6560
rect 31720 6496 31736 6560
rect 31800 6496 31808 6560
rect 31488 6495 31808 6496
rect 51850 6560 52170 6561
rect 51850 6496 51858 6560
rect 51922 6496 51938 6560
rect 52002 6496 52018 6560
rect 52082 6496 52098 6560
rect 52162 6496 52170 6560
rect 51850 6495 52170 6496
rect 20069 6490 20135 6493
rect 28533 6490 28599 6493
rect 20069 6488 28599 6490
rect 20069 6432 20074 6488
rect 20130 6432 28538 6488
rect 28594 6432 28599 6488
rect 20069 6430 28599 6432
rect 20069 6427 20135 6430
rect 28533 6427 28599 6430
rect 41689 6490 41755 6493
rect 45921 6490 45987 6493
rect 41689 6488 45987 6490
rect 41689 6432 41694 6488
rect 41750 6432 45926 6488
rect 45982 6432 45987 6488
rect 41689 6430 45987 6432
rect 41689 6427 41755 6430
rect 45921 6427 45987 6430
rect 51257 6490 51323 6493
rect 51257 6488 51642 6490
rect 51257 6432 51262 6488
rect 51318 6432 51642 6488
rect 51257 6430 51642 6432
rect 51257 6427 51323 6430
rect 20345 6354 20411 6357
rect 42149 6354 42215 6357
rect 20345 6352 42215 6354
rect 20345 6296 20350 6352
rect 20406 6296 42154 6352
rect 42210 6296 42215 6352
rect 20345 6294 42215 6296
rect 20345 6291 20411 6294
rect 42149 6291 42215 6294
rect 50705 6354 50771 6357
rect 51165 6354 51231 6357
rect 50705 6352 51231 6354
rect 50705 6296 50710 6352
rect 50766 6296 51170 6352
rect 51226 6296 51231 6352
rect 50705 6294 51231 6296
rect 51582 6354 51642 6430
rect 53741 6354 53807 6357
rect 51582 6352 53807 6354
rect 51582 6296 53746 6352
rect 53802 6296 53807 6352
rect 51582 6294 53807 6296
rect 50705 6291 50771 6294
rect 51165 6291 51231 6294
rect 53741 6291 53807 6294
rect 53925 6354 53991 6357
rect 55121 6354 55187 6357
rect 53925 6352 55187 6354
rect 53925 6296 53930 6352
rect 53986 6296 55126 6352
rect 55182 6296 55187 6352
rect 53925 6294 55187 6296
rect 53925 6291 53991 6294
rect 55121 6291 55187 6294
rect 2681 6218 2747 6221
rect 21725 6218 21791 6221
rect 2681 6216 21791 6218
rect 2681 6160 2686 6216
rect 2742 6160 21730 6216
rect 21786 6160 21791 6216
rect 2681 6158 21791 6160
rect 2681 6155 2747 6158
rect 21725 6155 21791 6158
rect 31201 6218 31267 6221
rect 32581 6218 32647 6221
rect 31201 6216 32647 6218
rect 31201 6160 31206 6216
rect 31262 6160 32586 6216
rect 32642 6160 32647 6216
rect 31201 6158 32647 6160
rect 31201 6155 31267 6158
rect 32581 6155 32647 6158
rect 49509 6218 49575 6221
rect 52269 6218 52335 6221
rect 49509 6216 52335 6218
rect 49509 6160 49514 6216
rect 49570 6160 52274 6216
rect 52330 6160 52335 6216
rect 49509 6158 52335 6160
rect 49509 6155 49575 6158
rect 52269 6155 52335 6158
rect 30281 6082 30347 6085
rect 31753 6082 31819 6085
rect 30281 6080 31819 6082
rect 30281 6024 30286 6080
rect 30342 6024 31758 6080
rect 31814 6024 31819 6080
rect 30281 6022 31819 6024
rect 30281 6019 30347 6022
rect 31753 6019 31819 6022
rect 49325 6082 49391 6085
rect 54661 6082 54727 6085
rect 49325 6080 54727 6082
rect 49325 6024 49330 6080
rect 49386 6024 54666 6080
rect 54722 6024 54727 6080
rect 49325 6022 54727 6024
rect 49325 6019 49391 6022
rect 54661 6019 54727 6022
rect 21306 6016 21626 6017
rect 21306 5952 21314 6016
rect 21378 5952 21394 6016
rect 21458 5952 21474 6016
rect 21538 5952 21554 6016
rect 21618 5952 21626 6016
rect 21306 5951 21626 5952
rect 41669 6016 41989 6017
rect 41669 5952 41677 6016
rect 41741 5952 41757 6016
rect 41821 5952 41837 6016
rect 41901 5952 41917 6016
rect 41981 5952 41989 6016
rect 41669 5951 41989 5952
rect 27153 5946 27219 5949
rect 31293 5946 31359 5949
rect 27153 5944 31359 5946
rect 27153 5888 27158 5944
rect 27214 5888 31298 5944
rect 31354 5888 31359 5944
rect 27153 5886 31359 5888
rect 27153 5883 27219 5886
rect 31293 5883 31359 5886
rect 49417 5946 49483 5949
rect 53557 5946 53623 5949
rect 49417 5944 53623 5946
rect 49417 5888 49422 5944
rect 49478 5888 53562 5944
rect 53618 5888 53623 5944
rect 49417 5886 53623 5888
rect 49417 5883 49483 5886
rect 53557 5883 53623 5886
rect 30925 5810 30991 5813
rect 32397 5810 32463 5813
rect 30925 5808 32463 5810
rect 30925 5752 30930 5808
rect 30986 5752 32402 5808
rect 32458 5752 32463 5808
rect 30925 5750 32463 5752
rect 30925 5747 30991 5750
rect 32397 5747 32463 5750
rect 45185 5810 45251 5813
rect 45645 5810 45711 5813
rect 45185 5808 45711 5810
rect 45185 5752 45190 5808
rect 45246 5752 45650 5808
rect 45706 5752 45711 5808
rect 45185 5750 45711 5752
rect 45185 5747 45251 5750
rect 45645 5747 45711 5750
rect 49233 5810 49299 5813
rect 52177 5810 52243 5813
rect 49233 5808 52243 5810
rect 49233 5752 49238 5808
rect 49294 5752 52182 5808
rect 52238 5752 52243 5808
rect 49233 5750 52243 5752
rect 49233 5747 49299 5750
rect 52177 5747 52243 5750
rect 30557 5674 30623 5677
rect 31845 5674 31911 5677
rect 30557 5672 31911 5674
rect 30557 5616 30562 5672
rect 30618 5616 31850 5672
rect 31906 5616 31911 5672
rect 30557 5614 31911 5616
rect 30557 5611 30623 5614
rect 31845 5611 31911 5614
rect 0 5538 800 5568
rect 2773 5538 2839 5541
rect 0 5536 2839 5538
rect 0 5480 2778 5536
rect 2834 5480 2839 5536
rect 0 5478 2839 5480
rect 0 5448 800 5478
rect 2773 5475 2839 5478
rect 21173 5538 21239 5541
rect 28257 5538 28323 5541
rect 21173 5536 28323 5538
rect 21173 5480 21178 5536
rect 21234 5480 28262 5536
rect 28318 5480 28323 5536
rect 21173 5478 28323 5480
rect 21173 5475 21239 5478
rect 28257 5475 28323 5478
rect 28809 5538 28875 5541
rect 29361 5538 29427 5541
rect 28809 5536 29427 5538
rect 28809 5480 28814 5536
rect 28870 5480 29366 5536
rect 29422 5480 29427 5536
rect 28809 5478 29427 5480
rect 28809 5475 28875 5478
rect 29361 5475 29427 5478
rect 37222 5476 37228 5540
rect 37292 5538 37298 5540
rect 46749 5538 46815 5541
rect 37292 5536 46815 5538
rect 37292 5480 46754 5536
rect 46810 5480 46815 5536
rect 37292 5478 46815 5480
rect 37292 5476 37298 5478
rect 46749 5475 46815 5478
rect 11125 5472 11445 5473
rect 11125 5408 11133 5472
rect 11197 5408 11213 5472
rect 11277 5408 11293 5472
rect 11357 5408 11373 5472
rect 11437 5408 11445 5472
rect 11125 5407 11445 5408
rect 31488 5472 31808 5473
rect 31488 5408 31496 5472
rect 31560 5408 31576 5472
rect 31640 5408 31656 5472
rect 31720 5408 31736 5472
rect 31800 5408 31808 5472
rect 31488 5407 31808 5408
rect 51850 5472 52170 5473
rect 51850 5408 51858 5472
rect 51922 5408 51938 5472
rect 52002 5408 52018 5472
rect 52082 5408 52098 5472
rect 52162 5408 52170 5472
rect 51850 5407 52170 5408
rect 7833 5266 7899 5269
rect 13445 5266 13511 5269
rect 7833 5264 13511 5266
rect 7833 5208 7838 5264
rect 7894 5208 13450 5264
rect 13506 5208 13511 5264
rect 7833 5206 13511 5208
rect 7833 5203 7899 5206
rect 13445 5203 13511 5206
rect 24025 5266 24091 5269
rect 41413 5266 41479 5269
rect 47485 5266 47551 5269
rect 24025 5264 29010 5266
rect 24025 5208 24030 5264
rect 24086 5232 29010 5264
rect 41413 5264 47551 5266
rect 24086 5208 29194 5232
rect 24025 5206 29194 5208
rect 24025 5203 24091 5206
rect 28950 5172 29194 5206
rect 41413 5208 41418 5264
rect 41474 5208 47490 5264
rect 47546 5208 47551 5264
rect 41413 5206 47551 5208
rect 41413 5203 41479 5206
rect 47485 5203 47551 5206
rect 10961 5130 11027 5133
rect 25497 5130 25563 5133
rect 10961 5128 25563 5130
rect 10961 5072 10966 5128
rect 11022 5072 25502 5128
rect 25558 5072 25563 5128
rect 10961 5070 25563 5072
rect 29134 5130 29194 5172
rect 37222 5130 37228 5132
rect 29134 5070 37228 5130
rect 10961 5067 11027 5070
rect 25497 5067 25563 5070
rect 37222 5068 37228 5070
rect 37292 5068 37298 5132
rect 46749 5130 46815 5133
rect 46933 5130 46999 5133
rect 46749 5128 46999 5130
rect 46749 5072 46754 5128
rect 46810 5072 46938 5128
rect 46994 5072 46999 5128
rect 46749 5070 46999 5072
rect 46749 5067 46815 5070
rect 46933 5067 46999 5070
rect 21306 4928 21626 4929
rect 21306 4864 21314 4928
rect 21378 4864 21394 4928
rect 21458 4864 21474 4928
rect 21538 4864 21554 4928
rect 21618 4864 21626 4928
rect 21306 4863 21626 4864
rect 41669 4928 41989 4929
rect 41669 4864 41677 4928
rect 41741 4864 41757 4928
rect 41821 4864 41837 4928
rect 41901 4864 41917 4928
rect 41981 4864 41989 4928
rect 41669 4863 41989 4864
rect 30189 4858 30255 4861
rect 32489 4858 32555 4861
rect 30189 4856 32555 4858
rect 30189 4800 30194 4856
rect 30250 4800 32494 4856
rect 32550 4800 32555 4856
rect 30189 4798 32555 4800
rect 30189 4795 30255 4798
rect 32489 4795 32555 4798
rect 5809 4722 5875 4725
rect 12801 4722 12867 4725
rect 5809 4720 12867 4722
rect 5809 4664 5814 4720
rect 5870 4664 12806 4720
rect 12862 4664 12867 4720
rect 5809 4662 12867 4664
rect 5809 4659 5875 4662
rect 12801 4659 12867 4662
rect 12157 4586 12223 4589
rect 18781 4586 18847 4589
rect 18965 4586 19031 4589
rect 12157 4584 19031 4586
rect 12157 4528 12162 4584
rect 12218 4528 18786 4584
rect 18842 4528 18970 4584
rect 19026 4528 19031 4584
rect 12157 4526 19031 4528
rect 12157 4523 12223 4526
rect 18781 4523 18847 4526
rect 18965 4523 19031 4526
rect 31017 4586 31083 4589
rect 35341 4586 35407 4589
rect 31017 4584 35407 4586
rect 31017 4528 31022 4584
rect 31078 4528 35346 4584
rect 35402 4528 35407 4584
rect 31017 4526 35407 4528
rect 31017 4523 31083 4526
rect 35341 4523 35407 4526
rect 11125 4384 11445 4385
rect 11125 4320 11133 4384
rect 11197 4320 11213 4384
rect 11277 4320 11293 4384
rect 11357 4320 11373 4384
rect 11437 4320 11445 4384
rect 11125 4319 11445 4320
rect 31488 4384 31808 4385
rect 31488 4320 31496 4384
rect 31560 4320 31576 4384
rect 31640 4320 31656 4384
rect 31720 4320 31736 4384
rect 31800 4320 31808 4384
rect 31488 4319 31808 4320
rect 51850 4384 52170 4385
rect 51850 4320 51858 4384
rect 51922 4320 51938 4384
rect 52002 4320 52018 4384
rect 52082 4320 52098 4384
rect 52162 4320 52170 4384
rect 51850 4319 52170 4320
rect 18229 4314 18295 4317
rect 19241 4314 19307 4317
rect 18229 4312 19307 4314
rect 18229 4256 18234 4312
rect 18290 4256 19246 4312
rect 19302 4256 19307 4312
rect 18229 4254 19307 4256
rect 18229 4251 18295 4254
rect 19241 4251 19307 4254
rect 9949 4178 10015 4181
rect 10685 4178 10751 4181
rect 19333 4178 19399 4181
rect 23933 4178 23999 4181
rect 32949 4178 33015 4181
rect 9949 4176 23999 4178
rect 9949 4120 9954 4176
rect 10010 4120 10690 4176
rect 10746 4120 19338 4176
rect 19394 4120 23938 4176
rect 23994 4120 23999 4176
rect 9949 4118 23999 4120
rect 9949 4115 10015 4118
rect 10685 4115 10751 4118
rect 19333 4115 19399 4118
rect 23933 4115 23999 4118
rect 30422 4176 33015 4178
rect 30422 4120 32954 4176
rect 33010 4120 33015 4176
rect 30422 4118 33015 4120
rect 4061 4042 4127 4045
rect 20529 4042 20595 4045
rect 4061 4040 20595 4042
rect 4061 3984 4066 4040
rect 4122 3984 20534 4040
rect 20590 3984 20595 4040
rect 4061 3982 20595 3984
rect 4061 3979 4127 3982
rect 20529 3979 20595 3982
rect 22921 4042 22987 4045
rect 30422 4042 30482 4118
rect 32949 4115 33015 4118
rect 22921 4040 30482 4042
rect 22921 3984 22926 4040
rect 22982 3984 30482 4040
rect 22921 3982 30482 3984
rect 30649 4042 30715 4045
rect 56501 4042 56567 4045
rect 30649 4040 56567 4042
rect 30649 3984 30654 4040
rect 30710 3984 56506 4040
rect 56562 3984 56567 4040
rect 30649 3982 56567 3984
rect 22921 3979 22987 3982
rect 30649 3979 30715 3982
rect 56501 3979 56567 3982
rect 15285 3906 15351 3909
rect 19149 3906 19215 3909
rect 15285 3904 19215 3906
rect 15285 3848 15290 3904
rect 15346 3848 19154 3904
rect 19210 3848 19215 3904
rect 15285 3846 19215 3848
rect 15285 3843 15351 3846
rect 19149 3843 19215 3846
rect 26785 3906 26851 3909
rect 36813 3906 36879 3909
rect 26785 3904 36879 3906
rect 26785 3848 26790 3904
rect 26846 3848 36818 3904
rect 36874 3848 36879 3904
rect 26785 3846 36879 3848
rect 26785 3843 26851 3846
rect 36813 3843 36879 3846
rect 21306 3840 21626 3841
rect 21306 3776 21314 3840
rect 21378 3776 21394 3840
rect 21458 3776 21474 3840
rect 21538 3776 21554 3840
rect 21618 3776 21626 3840
rect 21306 3775 21626 3776
rect 41669 3840 41989 3841
rect 41669 3776 41677 3840
rect 41741 3776 41757 3840
rect 41821 3776 41837 3840
rect 41901 3776 41917 3840
rect 41981 3776 41989 3840
rect 41669 3775 41989 3776
rect 1209 3770 1275 3773
rect 9765 3770 9831 3773
rect 1209 3768 9831 3770
rect 1209 3712 1214 3768
rect 1270 3712 9770 3768
rect 9826 3712 9831 3768
rect 1209 3710 9831 3712
rect 1209 3707 1275 3710
rect 9765 3707 9831 3710
rect 24577 3770 24643 3773
rect 31661 3770 31727 3773
rect 24577 3768 31727 3770
rect 24577 3712 24582 3768
rect 24638 3712 31666 3768
rect 31722 3712 31727 3768
rect 24577 3710 31727 3712
rect 24577 3707 24643 3710
rect 31661 3707 31727 3710
rect 31845 3770 31911 3773
rect 36261 3770 36327 3773
rect 31845 3768 36327 3770
rect 31845 3712 31850 3768
rect 31906 3712 36266 3768
rect 36322 3712 36327 3768
rect 31845 3710 36327 3712
rect 31845 3707 31911 3710
rect 36261 3707 36327 3710
rect 6361 3634 6427 3637
rect 26969 3634 27035 3637
rect 6361 3632 27035 3634
rect 6361 3576 6366 3632
rect 6422 3576 26974 3632
rect 27030 3576 27035 3632
rect 6361 3574 27035 3576
rect 6361 3571 6427 3574
rect 26969 3571 27035 3574
rect 27337 3634 27403 3637
rect 34697 3634 34763 3637
rect 27337 3632 34763 3634
rect 27337 3576 27342 3632
rect 27398 3576 34702 3632
rect 34758 3576 34763 3632
rect 27337 3574 34763 3576
rect 27337 3571 27403 3574
rect 34697 3571 34763 3574
rect 34973 3634 35039 3637
rect 53097 3634 53163 3637
rect 34973 3632 53163 3634
rect 34973 3576 34978 3632
rect 35034 3576 53102 3632
rect 53158 3576 53163 3632
rect 34973 3574 53163 3576
rect 34973 3571 35039 3574
rect 53097 3571 53163 3574
rect 54017 3634 54083 3637
rect 56869 3634 56935 3637
rect 54017 3632 56935 3634
rect 54017 3576 54022 3632
rect 54078 3576 56874 3632
rect 56930 3576 56935 3632
rect 54017 3574 56935 3576
rect 54017 3571 54083 3574
rect 56869 3571 56935 3574
rect 3785 3498 3851 3501
rect 35525 3498 35591 3501
rect 3785 3496 35591 3498
rect 3785 3440 3790 3496
rect 3846 3440 35530 3496
rect 35586 3440 35591 3496
rect 3785 3438 35591 3440
rect 3785 3435 3851 3438
rect 35525 3435 35591 3438
rect 39021 3498 39087 3501
rect 42057 3498 42123 3501
rect 39021 3496 42123 3498
rect 39021 3440 39026 3496
rect 39082 3440 42062 3496
rect 42118 3440 42123 3496
rect 39021 3438 42123 3440
rect 39021 3435 39087 3438
rect 42057 3435 42123 3438
rect 0 3362 800 3392
rect 4061 3362 4127 3365
rect 0 3360 4127 3362
rect 0 3304 4066 3360
rect 4122 3304 4127 3360
rect 0 3302 4127 3304
rect 0 3272 800 3302
rect 4061 3299 4127 3302
rect 14733 3362 14799 3365
rect 17217 3362 17283 3365
rect 14733 3360 17283 3362
rect 14733 3304 14738 3360
rect 14794 3304 17222 3360
rect 17278 3304 17283 3360
rect 14733 3302 17283 3304
rect 14733 3299 14799 3302
rect 17217 3299 17283 3302
rect 22001 3362 22067 3365
rect 26785 3362 26851 3365
rect 22001 3360 26851 3362
rect 22001 3304 22006 3360
rect 22062 3304 26790 3360
rect 26846 3304 26851 3360
rect 22001 3302 26851 3304
rect 22001 3299 22067 3302
rect 26785 3299 26851 3302
rect 31937 3362 32003 3365
rect 34513 3362 34579 3365
rect 31937 3360 34579 3362
rect 31937 3304 31942 3360
rect 31998 3304 34518 3360
rect 34574 3304 34579 3360
rect 31937 3302 34579 3304
rect 31937 3299 32003 3302
rect 34513 3299 34579 3302
rect 34697 3362 34763 3365
rect 41321 3362 41387 3365
rect 34697 3360 41387 3362
rect 34697 3304 34702 3360
rect 34758 3304 41326 3360
rect 41382 3304 41387 3360
rect 34697 3302 41387 3304
rect 34697 3299 34763 3302
rect 41321 3299 41387 3302
rect 11125 3296 11445 3297
rect 11125 3232 11133 3296
rect 11197 3232 11213 3296
rect 11277 3232 11293 3296
rect 11357 3232 11373 3296
rect 11437 3232 11445 3296
rect 11125 3231 11445 3232
rect 31488 3296 31808 3297
rect 31488 3232 31496 3296
rect 31560 3232 31576 3296
rect 31640 3232 31656 3296
rect 31720 3232 31736 3296
rect 31800 3232 31808 3296
rect 31488 3231 31808 3232
rect 51850 3296 52170 3297
rect 51850 3232 51858 3296
rect 51922 3232 51938 3296
rect 52002 3232 52018 3296
rect 52082 3232 52098 3296
rect 52162 3232 52170 3296
rect 51850 3231 52170 3232
rect 23749 3226 23815 3229
rect 31293 3226 31359 3229
rect 23749 3224 31359 3226
rect 23749 3168 23754 3224
rect 23810 3168 31298 3224
rect 31354 3168 31359 3224
rect 23749 3166 31359 3168
rect 23749 3163 23815 3166
rect 31293 3163 31359 3166
rect 34237 3226 34303 3229
rect 48681 3226 48747 3229
rect 34237 3224 48747 3226
rect 34237 3168 34242 3224
rect 34298 3168 48686 3224
rect 48742 3168 48747 3224
rect 34237 3166 48747 3168
rect 34237 3163 34303 3166
rect 48681 3163 48747 3166
rect 4705 3090 4771 3093
rect 22553 3090 22619 3093
rect 4705 3088 22619 3090
rect 4705 3032 4710 3088
rect 4766 3032 22558 3088
rect 22614 3032 22619 3088
rect 4705 3030 22619 3032
rect 4705 3027 4771 3030
rect 22553 3027 22619 3030
rect 29821 3090 29887 3093
rect 55581 3090 55647 3093
rect 29821 3088 55647 3090
rect 29821 3032 29826 3088
rect 29882 3032 55586 3088
rect 55642 3032 55647 3088
rect 29821 3030 55647 3032
rect 29821 3027 29887 3030
rect 55581 3027 55647 3030
rect 5625 2954 5691 2957
rect 22369 2954 22435 2957
rect 5625 2952 22435 2954
rect 5625 2896 5630 2952
rect 5686 2896 22374 2952
rect 22430 2896 22435 2952
rect 5625 2894 22435 2896
rect 5625 2891 5691 2894
rect 22369 2891 22435 2894
rect 26325 2954 26391 2957
rect 38745 2954 38811 2957
rect 26325 2952 38811 2954
rect 26325 2896 26330 2952
rect 26386 2896 38750 2952
rect 38806 2896 38811 2952
rect 26325 2894 38811 2896
rect 26325 2891 26391 2894
rect 38745 2891 38811 2894
rect 52453 2954 52519 2957
rect 55581 2954 55647 2957
rect 52453 2952 55647 2954
rect 52453 2896 52458 2952
rect 52514 2896 55586 2952
rect 55642 2896 55647 2952
rect 52453 2894 55647 2896
rect 52453 2891 52519 2894
rect 55581 2891 55647 2894
rect 16757 2818 16823 2821
rect 18689 2818 18755 2821
rect 16757 2816 18755 2818
rect 16757 2760 16762 2816
rect 16818 2760 18694 2816
rect 18750 2760 18755 2816
rect 16757 2758 18755 2760
rect 16757 2755 16823 2758
rect 18689 2755 18755 2758
rect 26969 2818 27035 2821
rect 32305 2818 32371 2821
rect 26969 2816 32371 2818
rect 26969 2760 26974 2816
rect 27030 2760 32310 2816
rect 32366 2760 32371 2816
rect 26969 2758 32371 2760
rect 26969 2755 27035 2758
rect 32305 2755 32371 2758
rect 34513 2818 34579 2821
rect 36537 2818 36603 2821
rect 34513 2816 36603 2818
rect 34513 2760 34518 2816
rect 34574 2760 36542 2816
rect 36598 2760 36603 2816
rect 34513 2758 36603 2760
rect 34513 2755 34579 2758
rect 36537 2755 36603 2758
rect 21306 2752 21626 2753
rect 21306 2688 21314 2752
rect 21378 2688 21394 2752
rect 21458 2688 21474 2752
rect 21538 2688 21554 2752
rect 21618 2688 21626 2752
rect 21306 2687 21626 2688
rect 41669 2752 41989 2753
rect 41669 2688 41677 2752
rect 41741 2688 41757 2752
rect 41821 2688 41837 2752
rect 41901 2688 41917 2752
rect 41981 2688 41989 2752
rect 41669 2687 41989 2688
rect 16573 2682 16639 2685
rect 18781 2682 18847 2685
rect 16573 2680 18847 2682
rect 16573 2624 16578 2680
rect 16634 2624 18786 2680
rect 18842 2624 18847 2680
rect 16573 2622 18847 2624
rect 16573 2619 16639 2622
rect 18781 2619 18847 2622
rect 24117 2682 24183 2685
rect 30373 2682 30439 2685
rect 24117 2680 30439 2682
rect 24117 2624 24122 2680
rect 24178 2624 30378 2680
rect 30434 2624 30439 2680
rect 24117 2622 30439 2624
rect 24117 2619 24183 2622
rect 30373 2619 30439 2622
rect 33961 2682 34027 2685
rect 36169 2682 36235 2685
rect 33961 2680 36235 2682
rect 33961 2624 33966 2680
rect 34022 2624 36174 2680
rect 36230 2624 36235 2680
rect 33961 2622 36235 2624
rect 33961 2619 34027 2622
rect 36169 2619 36235 2622
rect 11125 2208 11445 2209
rect 11125 2144 11133 2208
rect 11197 2144 11213 2208
rect 11277 2144 11293 2208
rect 11357 2144 11373 2208
rect 11437 2144 11445 2208
rect 11125 2143 11445 2144
rect 31488 2208 31808 2209
rect 31488 2144 31496 2208
rect 31560 2144 31576 2208
rect 31640 2144 31656 2208
rect 31720 2144 31736 2208
rect 31800 2144 31808 2208
rect 31488 2143 31808 2144
rect 51850 2208 52170 2209
rect 51850 2144 51858 2208
rect 51922 2144 51938 2208
rect 52002 2144 52018 2208
rect 52082 2144 52098 2208
rect 52162 2144 52170 2208
rect 51850 2143 52170 2144
rect 0 1186 800 1216
rect 3417 1186 3483 1189
rect 0 1184 3483 1186
rect 0 1128 3422 1184
rect 3478 1128 3483 1184
rect 0 1126 3483 1128
rect 0 1096 800 1126
rect 3417 1123 3483 1126
<< via3 >>
rect 11133 17436 11197 17440
rect 11133 17380 11137 17436
rect 11137 17380 11193 17436
rect 11193 17380 11197 17436
rect 11133 17376 11197 17380
rect 11213 17436 11277 17440
rect 11213 17380 11217 17436
rect 11217 17380 11273 17436
rect 11273 17380 11277 17436
rect 11213 17376 11277 17380
rect 11293 17436 11357 17440
rect 11293 17380 11297 17436
rect 11297 17380 11353 17436
rect 11353 17380 11357 17436
rect 11293 17376 11357 17380
rect 11373 17436 11437 17440
rect 11373 17380 11377 17436
rect 11377 17380 11433 17436
rect 11433 17380 11437 17436
rect 11373 17376 11437 17380
rect 31496 17436 31560 17440
rect 31496 17380 31500 17436
rect 31500 17380 31556 17436
rect 31556 17380 31560 17436
rect 31496 17376 31560 17380
rect 31576 17436 31640 17440
rect 31576 17380 31580 17436
rect 31580 17380 31636 17436
rect 31636 17380 31640 17436
rect 31576 17376 31640 17380
rect 31656 17436 31720 17440
rect 31656 17380 31660 17436
rect 31660 17380 31716 17436
rect 31716 17380 31720 17436
rect 31656 17376 31720 17380
rect 31736 17436 31800 17440
rect 31736 17380 31740 17436
rect 31740 17380 31796 17436
rect 31796 17380 31800 17436
rect 31736 17376 31800 17380
rect 51858 17436 51922 17440
rect 51858 17380 51862 17436
rect 51862 17380 51918 17436
rect 51918 17380 51922 17436
rect 51858 17376 51922 17380
rect 51938 17436 52002 17440
rect 51938 17380 51942 17436
rect 51942 17380 51998 17436
rect 51998 17380 52002 17436
rect 51938 17376 52002 17380
rect 52018 17436 52082 17440
rect 52018 17380 52022 17436
rect 52022 17380 52078 17436
rect 52078 17380 52082 17436
rect 52018 17376 52082 17380
rect 52098 17436 52162 17440
rect 52098 17380 52102 17436
rect 52102 17380 52158 17436
rect 52158 17380 52162 17436
rect 52098 17376 52162 17380
rect 21314 16892 21378 16896
rect 21314 16836 21318 16892
rect 21318 16836 21374 16892
rect 21374 16836 21378 16892
rect 21314 16832 21378 16836
rect 21394 16892 21458 16896
rect 21394 16836 21398 16892
rect 21398 16836 21454 16892
rect 21454 16836 21458 16892
rect 21394 16832 21458 16836
rect 21474 16892 21538 16896
rect 21474 16836 21478 16892
rect 21478 16836 21534 16892
rect 21534 16836 21538 16892
rect 21474 16832 21538 16836
rect 21554 16892 21618 16896
rect 21554 16836 21558 16892
rect 21558 16836 21614 16892
rect 21614 16836 21618 16892
rect 21554 16832 21618 16836
rect 41677 16892 41741 16896
rect 41677 16836 41681 16892
rect 41681 16836 41737 16892
rect 41737 16836 41741 16892
rect 41677 16832 41741 16836
rect 41757 16892 41821 16896
rect 41757 16836 41761 16892
rect 41761 16836 41817 16892
rect 41817 16836 41821 16892
rect 41757 16832 41821 16836
rect 41837 16892 41901 16896
rect 41837 16836 41841 16892
rect 41841 16836 41897 16892
rect 41897 16836 41901 16892
rect 41837 16832 41901 16836
rect 41917 16892 41981 16896
rect 41917 16836 41921 16892
rect 41921 16836 41977 16892
rect 41977 16836 41981 16892
rect 41917 16832 41981 16836
rect 11133 16348 11197 16352
rect 11133 16292 11137 16348
rect 11137 16292 11193 16348
rect 11193 16292 11197 16348
rect 11133 16288 11197 16292
rect 11213 16348 11277 16352
rect 11213 16292 11217 16348
rect 11217 16292 11273 16348
rect 11273 16292 11277 16348
rect 11213 16288 11277 16292
rect 11293 16348 11357 16352
rect 11293 16292 11297 16348
rect 11297 16292 11353 16348
rect 11353 16292 11357 16348
rect 11293 16288 11357 16292
rect 11373 16348 11437 16352
rect 11373 16292 11377 16348
rect 11377 16292 11433 16348
rect 11433 16292 11437 16348
rect 11373 16288 11437 16292
rect 31496 16348 31560 16352
rect 31496 16292 31500 16348
rect 31500 16292 31556 16348
rect 31556 16292 31560 16348
rect 31496 16288 31560 16292
rect 31576 16348 31640 16352
rect 31576 16292 31580 16348
rect 31580 16292 31636 16348
rect 31636 16292 31640 16348
rect 31576 16288 31640 16292
rect 31656 16348 31720 16352
rect 31656 16292 31660 16348
rect 31660 16292 31716 16348
rect 31716 16292 31720 16348
rect 31656 16288 31720 16292
rect 31736 16348 31800 16352
rect 31736 16292 31740 16348
rect 31740 16292 31796 16348
rect 31796 16292 31800 16348
rect 31736 16288 31800 16292
rect 51858 16348 51922 16352
rect 51858 16292 51862 16348
rect 51862 16292 51918 16348
rect 51918 16292 51922 16348
rect 51858 16288 51922 16292
rect 51938 16348 52002 16352
rect 51938 16292 51942 16348
rect 51942 16292 51998 16348
rect 51998 16292 52002 16348
rect 51938 16288 52002 16292
rect 52018 16348 52082 16352
rect 52018 16292 52022 16348
rect 52022 16292 52078 16348
rect 52078 16292 52082 16348
rect 52018 16288 52082 16292
rect 52098 16348 52162 16352
rect 52098 16292 52102 16348
rect 52102 16292 52158 16348
rect 52158 16292 52162 16348
rect 52098 16288 52162 16292
rect 21314 15804 21378 15808
rect 21314 15748 21318 15804
rect 21318 15748 21374 15804
rect 21374 15748 21378 15804
rect 21314 15744 21378 15748
rect 21394 15804 21458 15808
rect 21394 15748 21398 15804
rect 21398 15748 21454 15804
rect 21454 15748 21458 15804
rect 21394 15744 21458 15748
rect 21474 15804 21538 15808
rect 21474 15748 21478 15804
rect 21478 15748 21534 15804
rect 21534 15748 21538 15804
rect 21474 15744 21538 15748
rect 21554 15804 21618 15808
rect 21554 15748 21558 15804
rect 21558 15748 21614 15804
rect 21614 15748 21618 15804
rect 21554 15744 21618 15748
rect 41677 15804 41741 15808
rect 41677 15748 41681 15804
rect 41681 15748 41737 15804
rect 41737 15748 41741 15804
rect 41677 15744 41741 15748
rect 41757 15804 41821 15808
rect 41757 15748 41761 15804
rect 41761 15748 41817 15804
rect 41817 15748 41821 15804
rect 41757 15744 41821 15748
rect 41837 15804 41901 15808
rect 41837 15748 41841 15804
rect 41841 15748 41897 15804
rect 41897 15748 41901 15804
rect 41837 15744 41901 15748
rect 41917 15804 41981 15808
rect 41917 15748 41921 15804
rect 41921 15748 41977 15804
rect 41977 15748 41981 15804
rect 41917 15744 41981 15748
rect 11133 15260 11197 15264
rect 11133 15204 11137 15260
rect 11137 15204 11193 15260
rect 11193 15204 11197 15260
rect 11133 15200 11197 15204
rect 11213 15260 11277 15264
rect 11213 15204 11217 15260
rect 11217 15204 11273 15260
rect 11273 15204 11277 15260
rect 11213 15200 11277 15204
rect 11293 15260 11357 15264
rect 11293 15204 11297 15260
rect 11297 15204 11353 15260
rect 11353 15204 11357 15260
rect 11293 15200 11357 15204
rect 11373 15260 11437 15264
rect 11373 15204 11377 15260
rect 11377 15204 11433 15260
rect 11433 15204 11437 15260
rect 11373 15200 11437 15204
rect 31496 15260 31560 15264
rect 31496 15204 31500 15260
rect 31500 15204 31556 15260
rect 31556 15204 31560 15260
rect 31496 15200 31560 15204
rect 31576 15260 31640 15264
rect 31576 15204 31580 15260
rect 31580 15204 31636 15260
rect 31636 15204 31640 15260
rect 31576 15200 31640 15204
rect 31656 15260 31720 15264
rect 31656 15204 31660 15260
rect 31660 15204 31716 15260
rect 31716 15204 31720 15260
rect 31656 15200 31720 15204
rect 31736 15260 31800 15264
rect 31736 15204 31740 15260
rect 31740 15204 31796 15260
rect 31796 15204 31800 15260
rect 31736 15200 31800 15204
rect 51858 15260 51922 15264
rect 51858 15204 51862 15260
rect 51862 15204 51918 15260
rect 51918 15204 51922 15260
rect 51858 15200 51922 15204
rect 51938 15260 52002 15264
rect 51938 15204 51942 15260
rect 51942 15204 51998 15260
rect 51998 15204 52002 15260
rect 51938 15200 52002 15204
rect 52018 15260 52082 15264
rect 52018 15204 52022 15260
rect 52022 15204 52078 15260
rect 52078 15204 52082 15260
rect 52018 15200 52082 15204
rect 52098 15260 52162 15264
rect 52098 15204 52102 15260
rect 52102 15204 52158 15260
rect 52158 15204 52162 15260
rect 52098 15200 52162 15204
rect 21314 14716 21378 14720
rect 21314 14660 21318 14716
rect 21318 14660 21374 14716
rect 21374 14660 21378 14716
rect 21314 14656 21378 14660
rect 21394 14716 21458 14720
rect 21394 14660 21398 14716
rect 21398 14660 21454 14716
rect 21454 14660 21458 14716
rect 21394 14656 21458 14660
rect 21474 14716 21538 14720
rect 21474 14660 21478 14716
rect 21478 14660 21534 14716
rect 21534 14660 21538 14716
rect 21474 14656 21538 14660
rect 21554 14716 21618 14720
rect 21554 14660 21558 14716
rect 21558 14660 21614 14716
rect 21614 14660 21618 14716
rect 21554 14656 21618 14660
rect 41677 14716 41741 14720
rect 41677 14660 41681 14716
rect 41681 14660 41737 14716
rect 41737 14660 41741 14716
rect 41677 14656 41741 14660
rect 41757 14716 41821 14720
rect 41757 14660 41761 14716
rect 41761 14660 41817 14716
rect 41817 14660 41821 14716
rect 41757 14656 41821 14660
rect 41837 14716 41901 14720
rect 41837 14660 41841 14716
rect 41841 14660 41897 14716
rect 41897 14660 41901 14716
rect 41837 14656 41901 14660
rect 41917 14716 41981 14720
rect 41917 14660 41921 14716
rect 41921 14660 41977 14716
rect 41977 14660 41981 14716
rect 41917 14656 41981 14660
rect 11133 14172 11197 14176
rect 11133 14116 11137 14172
rect 11137 14116 11193 14172
rect 11193 14116 11197 14172
rect 11133 14112 11197 14116
rect 11213 14172 11277 14176
rect 11213 14116 11217 14172
rect 11217 14116 11273 14172
rect 11273 14116 11277 14172
rect 11213 14112 11277 14116
rect 11293 14172 11357 14176
rect 11293 14116 11297 14172
rect 11297 14116 11353 14172
rect 11353 14116 11357 14172
rect 11293 14112 11357 14116
rect 11373 14172 11437 14176
rect 11373 14116 11377 14172
rect 11377 14116 11433 14172
rect 11433 14116 11437 14172
rect 11373 14112 11437 14116
rect 31496 14172 31560 14176
rect 31496 14116 31500 14172
rect 31500 14116 31556 14172
rect 31556 14116 31560 14172
rect 31496 14112 31560 14116
rect 31576 14172 31640 14176
rect 31576 14116 31580 14172
rect 31580 14116 31636 14172
rect 31636 14116 31640 14172
rect 31576 14112 31640 14116
rect 31656 14172 31720 14176
rect 31656 14116 31660 14172
rect 31660 14116 31716 14172
rect 31716 14116 31720 14172
rect 31656 14112 31720 14116
rect 31736 14172 31800 14176
rect 31736 14116 31740 14172
rect 31740 14116 31796 14172
rect 31796 14116 31800 14172
rect 31736 14112 31800 14116
rect 51858 14172 51922 14176
rect 51858 14116 51862 14172
rect 51862 14116 51918 14172
rect 51918 14116 51922 14172
rect 51858 14112 51922 14116
rect 51938 14172 52002 14176
rect 51938 14116 51942 14172
rect 51942 14116 51998 14172
rect 51998 14116 52002 14172
rect 51938 14112 52002 14116
rect 52018 14172 52082 14176
rect 52018 14116 52022 14172
rect 52022 14116 52078 14172
rect 52078 14116 52082 14172
rect 52018 14112 52082 14116
rect 52098 14172 52162 14176
rect 52098 14116 52102 14172
rect 52102 14116 52158 14172
rect 52158 14116 52162 14172
rect 52098 14112 52162 14116
rect 21314 13628 21378 13632
rect 21314 13572 21318 13628
rect 21318 13572 21374 13628
rect 21374 13572 21378 13628
rect 21314 13568 21378 13572
rect 21394 13628 21458 13632
rect 21394 13572 21398 13628
rect 21398 13572 21454 13628
rect 21454 13572 21458 13628
rect 21394 13568 21458 13572
rect 21474 13628 21538 13632
rect 21474 13572 21478 13628
rect 21478 13572 21534 13628
rect 21534 13572 21538 13628
rect 21474 13568 21538 13572
rect 21554 13628 21618 13632
rect 21554 13572 21558 13628
rect 21558 13572 21614 13628
rect 21614 13572 21618 13628
rect 21554 13568 21618 13572
rect 41677 13628 41741 13632
rect 41677 13572 41681 13628
rect 41681 13572 41737 13628
rect 41737 13572 41741 13628
rect 41677 13568 41741 13572
rect 41757 13628 41821 13632
rect 41757 13572 41761 13628
rect 41761 13572 41817 13628
rect 41817 13572 41821 13628
rect 41757 13568 41821 13572
rect 41837 13628 41901 13632
rect 41837 13572 41841 13628
rect 41841 13572 41897 13628
rect 41897 13572 41901 13628
rect 41837 13568 41901 13572
rect 41917 13628 41981 13632
rect 41917 13572 41921 13628
rect 41921 13572 41977 13628
rect 41977 13572 41981 13628
rect 41917 13568 41981 13572
rect 11133 13084 11197 13088
rect 11133 13028 11137 13084
rect 11137 13028 11193 13084
rect 11193 13028 11197 13084
rect 11133 13024 11197 13028
rect 11213 13084 11277 13088
rect 11213 13028 11217 13084
rect 11217 13028 11273 13084
rect 11273 13028 11277 13084
rect 11213 13024 11277 13028
rect 11293 13084 11357 13088
rect 11293 13028 11297 13084
rect 11297 13028 11353 13084
rect 11353 13028 11357 13084
rect 11293 13024 11357 13028
rect 11373 13084 11437 13088
rect 11373 13028 11377 13084
rect 11377 13028 11433 13084
rect 11433 13028 11437 13084
rect 11373 13024 11437 13028
rect 31496 13084 31560 13088
rect 31496 13028 31500 13084
rect 31500 13028 31556 13084
rect 31556 13028 31560 13084
rect 31496 13024 31560 13028
rect 31576 13084 31640 13088
rect 31576 13028 31580 13084
rect 31580 13028 31636 13084
rect 31636 13028 31640 13084
rect 31576 13024 31640 13028
rect 31656 13084 31720 13088
rect 31656 13028 31660 13084
rect 31660 13028 31716 13084
rect 31716 13028 31720 13084
rect 31656 13024 31720 13028
rect 31736 13084 31800 13088
rect 31736 13028 31740 13084
rect 31740 13028 31796 13084
rect 31796 13028 31800 13084
rect 31736 13024 31800 13028
rect 51858 13084 51922 13088
rect 51858 13028 51862 13084
rect 51862 13028 51918 13084
rect 51918 13028 51922 13084
rect 51858 13024 51922 13028
rect 51938 13084 52002 13088
rect 51938 13028 51942 13084
rect 51942 13028 51998 13084
rect 51998 13028 52002 13084
rect 51938 13024 52002 13028
rect 52018 13084 52082 13088
rect 52018 13028 52022 13084
rect 52022 13028 52078 13084
rect 52078 13028 52082 13084
rect 52018 13024 52082 13028
rect 52098 13084 52162 13088
rect 52098 13028 52102 13084
rect 52102 13028 52158 13084
rect 52158 13028 52162 13084
rect 52098 13024 52162 13028
rect 21314 12540 21378 12544
rect 21314 12484 21318 12540
rect 21318 12484 21374 12540
rect 21374 12484 21378 12540
rect 21314 12480 21378 12484
rect 21394 12540 21458 12544
rect 21394 12484 21398 12540
rect 21398 12484 21454 12540
rect 21454 12484 21458 12540
rect 21394 12480 21458 12484
rect 21474 12540 21538 12544
rect 21474 12484 21478 12540
rect 21478 12484 21534 12540
rect 21534 12484 21538 12540
rect 21474 12480 21538 12484
rect 21554 12540 21618 12544
rect 21554 12484 21558 12540
rect 21558 12484 21614 12540
rect 21614 12484 21618 12540
rect 21554 12480 21618 12484
rect 41677 12540 41741 12544
rect 41677 12484 41681 12540
rect 41681 12484 41737 12540
rect 41737 12484 41741 12540
rect 41677 12480 41741 12484
rect 41757 12540 41821 12544
rect 41757 12484 41761 12540
rect 41761 12484 41817 12540
rect 41817 12484 41821 12540
rect 41757 12480 41821 12484
rect 41837 12540 41901 12544
rect 41837 12484 41841 12540
rect 41841 12484 41897 12540
rect 41897 12484 41901 12540
rect 41837 12480 41901 12484
rect 41917 12540 41981 12544
rect 41917 12484 41921 12540
rect 41921 12484 41977 12540
rect 41977 12484 41981 12540
rect 41917 12480 41981 12484
rect 11133 11996 11197 12000
rect 11133 11940 11137 11996
rect 11137 11940 11193 11996
rect 11193 11940 11197 11996
rect 11133 11936 11197 11940
rect 11213 11996 11277 12000
rect 11213 11940 11217 11996
rect 11217 11940 11273 11996
rect 11273 11940 11277 11996
rect 11213 11936 11277 11940
rect 11293 11996 11357 12000
rect 11293 11940 11297 11996
rect 11297 11940 11353 11996
rect 11353 11940 11357 11996
rect 11293 11936 11357 11940
rect 11373 11996 11437 12000
rect 11373 11940 11377 11996
rect 11377 11940 11433 11996
rect 11433 11940 11437 11996
rect 11373 11936 11437 11940
rect 31496 11996 31560 12000
rect 31496 11940 31500 11996
rect 31500 11940 31556 11996
rect 31556 11940 31560 11996
rect 31496 11936 31560 11940
rect 31576 11996 31640 12000
rect 31576 11940 31580 11996
rect 31580 11940 31636 11996
rect 31636 11940 31640 11996
rect 31576 11936 31640 11940
rect 31656 11996 31720 12000
rect 31656 11940 31660 11996
rect 31660 11940 31716 11996
rect 31716 11940 31720 11996
rect 31656 11936 31720 11940
rect 31736 11996 31800 12000
rect 31736 11940 31740 11996
rect 31740 11940 31796 11996
rect 31796 11940 31800 11996
rect 31736 11936 31800 11940
rect 51858 11996 51922 12000
rect 51858 11940 51862 11996
rect 51862 11940 51918 11996
rect 51918 11940 51922 11996
rect 51858 11936 51922 11940
rect 51938 11996 52002 12000
rect 51938 11940 51942 11996
rect 51942 11940 51998 11996
rect 51998 11940 52002 11996
rect 51938 11936 52002 11940
rect 52018 11996 52082 12000
rect 52018 11940 52022 11996
rect 52022 11940 52078 11996
rect 52078 11940 52082 11996
rect 52018 11936 52082 11940
rect 52098 11996 52162 12000
rect 52098 11940 52102 11996
rect 52102 11940 52158 11996
rect 52158 11940 52162 11996
rect 52098 11936 52162 11940
rect 21314 11452 21378 11456
rect 21314 11396 21318 11452
rect 21318 11396 21374 11452
rect 21374 11396 21378 11452
rect 21314 11392 21378 11396
rect 21394 11452 21458 11456
rect 21394 11396 21398 11452
rect 21398 11396 21454 11452
rect 21454 11396 21458 11452
rect 21394 11392 21458 11396
rect 21474 11452 21538 11456
rect 21474 11396 21478 11452
rect 21478 11396 21534 11452
rect 21534 11396 21538 11452
rect 21474 11392 21538 11396
rect 21554 11452 21618 11456
rect 21554 11396 21558 11452
rect 21558 11396 21614 11452
rect 21614 11396 21618 11452
rect 21554 11392 21618 11396
rect 41677 11452 41741 11456
rect 41677 11396 41681 11452
rect 41681 11396 41737 11452
rect 41737 11396 41741 11452
rect 41677 11392 41741 11396
rect 41757 11452 41821 11456
rect 41757 11396 41761 11452
rect 41761 11396 41817 11452
rect 41817 11396 41821 11452
rect 41757 11392 41821 11396
rect 41837 11452 41901 11456
rect 41837 11396 41841 11452
rect 41841 11396 41897 11452
rect 41897 11396 41901 11452
rect 41837 11392 41901 11396
rect 41917 11452 41981 11456
rect 41917 11396 41921 11452
rect 41921 11396 41977 11452
rect 41977 11396 41981 11452
rect 41917 11392 41981 11396
rect 11133 10908 11197 10912
rect 11133 10852 11137 10908
rect 11137 10852 11193 10908
rect 11193 10852 11197 10908
rect 11133 10848 11197 10852
rect 11213 10908 11277 10912
rect 11213 10852 11217 10908
rect 11217 10852 11273 10908
rect 11273 10852 11277 10908
rect 11213 10848 11277 10852
rect 11293 10908 11357 10912
rect 11293 10852 11297 10908
rect 11297 10852 11353 10908
rect 11353 10852 11357 10908
rect 11293 10848 11357 10852
rect 11373 10908 11437 10912
rect 11373 10852 11377 10908
rect 11377 10852 11433 10908
rect 11433 10852 11437 10908
rect 11373 10848 11437 10852
rect 31496 10908 31560 10912
rect 31496 10852 31500 10908
rect 31500 10852 31556 10908
rect 31556 10852 31560 10908
rect 31496 10848 31560 10852
rect 31576 10908 31640 10912
rect 31576 10852 31580 10908
rect 31580 10852 31636 10908
rect 31636 10852 31640 10908
rect 31576 10848 31640 10852
rect 31656 10908 31720 10912
rect 31656 10852 31660 10908
rect 31660 10852 31716 10908
rect 31716 10852 31720 10908
rect 31656 10848 31720 10852
rect 31736 10908 31800 10912
rect 31736 10852 31740 10908
rect 31740 10852 31796 10908
rect 31796 10852 31800 10908
rect 31736 10848 31800 10852
rect 51858 10908 51922 10912
rect 51858 10852 51862 10908
rect 51862 10852 51918 10908
rect 51918 10852 51922 10908
rect 51858 10848 51922 10852
rect 51938 10908 52002 10912
rect 51938 10852 51942 10908
rect 51942 10852 51998 10908
rect 51998 10852 52002 10908
rect 51938 10848 52002 10852
rect 52018 10908 52082 10912
rect 52018 10852 52022 10908
rect 52022 10852 52078 10908
rect 52078 10852 52082 10908
rect 52018 10848 52082 10852
rect 52098 10908 52162 10912
rect 52098 10852 52102 10908
rect 52102 10852 52158 10908
rect 52158 10852 52162 10908
rect 52098 10848 52162 10852
rect 21314 10364 21378 10368
rect 21314 10308 21318 10364
rect 21318 10308 21374 10364
rect 21374 10308 21378 10364
rect 21314 10304 21378 10308
rect 21394 10364 21458 10368
rect 21394 10308 21398 10364
rect 21398 10308 21454 10364
rect 21454 10308 21458 10364
rect 21394 10304 21458 10308
rect 21474 10364 21538 10368
rect 21474 10308 21478 10364
rect 21478 10308 21534 10364
rect 21534 10308 21538 10364
rect 21474 10304 21538 10308
rect 21554 10364 21618 10368
rect 21554 10308 21558 10364
rect 21558 10308 21614 10364
rect 21614 10308 21618 10364
rect 21554 10304 21618 10308
rect 41677 10364 41741 10368
rect 41677 10308 41681 10364
rect 41681 10308 41737 10364
rect 41737 10308 41741 10364
rect 41677 10304 41741 10308
rect 41757 10364 41821 10368
rect 41757 10308 41761 10364
rect 41761 10308 41817 10364
rect 41817 10308 41821 10364
rect 41757 10304 41821 10308
rect 41837 10364 41901 10368
rect 41837 10308 41841 10364
rect 41841 10308 41897 10364
rect 41897 10308 41901 10364
rect 41837 10304 41901 10308
rect 41917 10364 41981 10368
rect 41917 10308 41921 10364
rect 41921 10308 41977 10364
rect 41977 10308 41981 10364
rect 41917 10304 41981 10308
rect 11133 9820 11197 9824
rect 11133 9764 11137 9820
rect 11137 9764 11193 9820
rect 11193 9764 11197 9820
rect 11133 9760 11197 9764
rect 11213 9820 11277 9824
rect 11213 9764 11217 9820
rect 11217 9764 11273 9820
rect 11273 9764 11277 9820
rect 11213 9760 11277 9764
rect 11293 9820 11357 9824
rect 11293 9764 11297 9820
rect 11297 9764 11353 9820
rect 11353 9764 11357 9820
rect 11293 9760 11357 9764
rect 11373 9820 11437 9824
rect 11373 9764 11377 9820
rect 11377 9764 11433 9820
rect 11433 9764 11437 9820
rect 11373 9760 11437 9764
rect 31496 9820 31560 9824
rect 31496 9764 31500 9820
rect 31500 9764 31556 9820
rect 31556 9764 31560 9820
rect 31496 9760 31560 9764
rect 31576 9820 31640 9824
rect 31576 9764 31580 9820
rect 31580 9764 31636 9820
rect 31636 9764 31640 9820
rect 31576 9760 31640 9764
rect 31656 9820 31720 9824
rect 31656 9764 31660 9820
rect 31660 9764 31716 9820
rect 31716 9764 31720 9820
rect 31656 9760 31720 9764
rect 31736 9820 31800 9824
rect 31736 9764 31740 9820
rect 31740 9764 31796 9820
rect 31796 9764 31800 9820
rect 31736 9760 31800 9764
rect 51858 9820 51922 9824
rect 51858 9764 51862 9820
rect 51862 9764 51918 9820
rect 51918 9764 51922 9820
rect 51858 9760 51922 9764
rect 51938 9820 52002 9824
rect 51938 9764 51942 9820
rect 51942 9764 51998 9820
rect 51998 9764 52002 9820
rect 51938 9760 52002 9764
rect 52018 9820 52082 9824
rect 52018 9764 52022 9820
rect 52022 9764 52078 9820
rect 52078 9764 52082 9820
rect 52018 9760 52082 9764
rect 52098 9820 52162 9824
rect 52098 9764 52102 9820
rect 52102 9764 52158 9820
rect 52158 9764 52162 9820
rect 52098 9760 52162 9764
rect 21314 9276 21378 9280
rect 21314 9220 21318 9276
rect 21318 9220 21374 9276
rect 21374 9220 21378 9276
rect 21314 9216 21378 9220
rect 21394 9276 21458 9280
rect 21394 9220 21398 9276
rect 21398 9220 21454 9276
rect 21454 9220 21458 9276
rect 21394 9216 21458 9220
rect 21474 9276 21538 9280
rect 21474 9220 21478 9276
rect 21478 9220 21534 9276
rect 21534 9220 21538 9276
rect 21474 9216 21538 9220
rect 21554 9276 21618 9280
rect 21554 9220 21558 9276
rect 21558 9220 21614 9276
rect 21614 9220 21618 9276
rect 21554 9216 21618 9220
rect 41677 9276 41741 9280
rect 41677 9220 41681 9276
rect 41681 9220 41737 9276
rect 41737 9220 41741 9276
rect 41677 9216 41741 9220
rect 41757 9276 41821 9280
rect 41757 9220 41761 9276
rect 41761 9220 41817 9276
rect 41817 9220 41821 9276
rect 41757 9216 41821 9220
rect 41837 9276 41901 9280
rect 41837 9220 41841 9276
rect 41841 9220 41897 9276
rect 41897 9220 41901 9276
rect 41837 9216 41901 9220
rect 41917 9276 41981 9280
rect 41917 9220 41921 9276
rect 41921 9220 41977 9276
rect 41977 9220 41981 9276
rect 41917 9216 41981 9220
rect 11133 8732 11197 8736
rect 11133 8676 11137 8732
rect 11137 8676 11193 8732
rect 11193 8676 11197 8732
rect 11133 8672 11197 8676
rect 11213 8732 11277 8736
rect 11213 8676 11217 8732
rect 11217 8676 11273 8732
rect 11273 8676 11277 8732
rect 11213 8672 11277 8676
rect 11293 8732 11357 8736
rect 11293 8676 11297 8732
rect 11297 8676 11353 8732
rect 11353 8676 11357 8732
rect 11293 8672 11357 8676
rect 11373 8732 11437 8736
rect 11373 8676 11377 8732
rect 11377 8676 11433 8732
rect 11433 8676 11437 8732
rect 11373 8672 11437 8676
rect 31496 8732 31560 8736
rect 31496 8676 31500 8732
rect 31500 8676 31556 8732
rect 31556 8676 31560 8732
rect 31496 8672 31560 8676
rect 31576 8732 31640 8736
rect 31576 8676 31580 8732
rect 31580 8676 31636 8732
rect 31636 8676 31640 8732
rect 31576 8672 31640 8676
rect 31656 8732 31720 8736
rect 31656 8676 31660 8732
rect 31660 8676 31716 8732
rect 31716 8676 31720 8732
rect 31656 8672 31720 8676
rect 31736 8732 31800 8736
rect 31736 8676 31740 8732
rect 31740 8676 31796 8732
rect 31796 8676 31800 8732
rect 31736 8672 31800 8676
rect 51858 8732 51922 8736
rect 51858 8676 51862 8732
rect 51862 8676 51918 8732
rect 51918 8676 51922 8732
rect 51858 8672 51922 8676
rect 51938 8732 52002 8736
rect 51938 8676 51942 8732
rect 51942 8676 51998 8732
rect 51998 8676 52002 8732
rect 51938 8672 52002 8676
rect 52018 8732 52082 8736
rect 52018 8676 52022 8732
rect 52022 8676 52078 8732
rect 52078 8676 52082 8732
rect 52018 8672 52082 8676
rect 52098 8732 52162 8736
rect 52098 8676 52102 8732
rect 52102 8676 52158 8732
rect 52158 8676 52162 8732
rect 52098 8672 52162 8676
rect 21314 8188 21378 8192
rect 21314 8132 21318 8188
rect 21318 8132 21374 8188
rect 21374 8132 21378 8188
rect 21314 8128 21378 8132
rect 21394 8188 21458 8192
rect 21394 8132 21398 8188
rect 21398 8132 21454 8188
rect 21454 8132 21458 8188
rect 21394 8128 21458 8132
rect 21474 8188 21538 8192
rect 21474 8132 21478 8188
rect 21478 8132 21534 8188
rect 21534 8132 21538 8188
rect 21474 8128 21538 8132
rect 21554 8188 21618 8192
rect 21554 8132 21558 8188
rect 21558 8132 21614 8188
rect 21614 8132 21618 8188
rect 21554 8128 21618 8132
rect 41677 8188 41741 8192
rect 41677 8132 41681 8188
rect 41681 8132 41737 8188
rect 41737 8132 41741 8188
rect 41677 8128 41741 8132
rect 41757 8188 41821 8192
rect 41757 8132 41761 8188
rect 41761 8132 41817 8188
rect 41817 8132 41821 8188
rect 41757 8128 41821 8132
rect 41837 8188 41901 8192
rect 41837 8132 41841 8188
rect 41841 8132 41897 8188
rect 41897 8132 41901 8188
rect 41837 8128 41901 8132
rect 41917 8188 41981 8192
rect 41917 8132 41921 8188
rect 41921 8132 41977 8188
rect 41977 8132 41981 8188
rect 41917 8128 41981 8132
rect 11133 7644 11197 7648
rect 11133 7588 11137 7644
rect 11137 7588 11193 7644
rect 11193 7588 11197 7644
rect 11133 7584 11197 7588
rect 11213 7644 11277 7648
rect 11213 7588 11217 7644
rect 11217 7588 11273 7644
rect 11273 7588 11277 7644
rect 11213 7584 11277 7588
rect 11293 7644 11357 7648
rect 11293 7588 11297 7644
rect 11297 7588 11353 7644
rect 11353 7588 11357 7644
rect 11293 7584 11357 7588
rect 11373 7644 11437 7648
rect 11373 7588 11377 7644
rect 11377 7588 11433 7644
rect 11433 7588 11437 7644
rect 11373 7584 11437 7588
rect 31496 7644 31560 7648
rect 31496 7588 31500 7644
rect 31500 7588 31556 7644
rect 31556 7588 31560 7644
rect 31496 7584 31560 7588
rect 31576 7644 31640 7648
rect 31576 7588 31580 7644
rect 31580 7588 31636 7644
rect 31636 7588 31640 7644
rect 31576 7584 31640 7588
rect 31656 7644 31720 7648
rect 31656 7588 31660 7644
rect 31660 7588 31716 7644
rect 31716 7588 31720 7644
rect 31656 7584 31720 7588
rect 31736 7644 31800 7648
rect 31736 7588 31740 7644
rect 31740 7588 31796 7644
rect 31796 7588 31800 7644
rect 31736 7584 31800 7588
rect 51858 7644 51922 7648
rect 51858 7588 51862 7644
rect 51862 7588 51918 7644
rect 51918 7588 51922 7644
rect 51858 7584 51922 7588
rect 51938 7644 52002 7648
rect 51938 7588 51942 7644
rect 51942 7588 51998 7644
rect 51998 7588 52002 7644
rect 51938 7584 52002 7588
rect 52018 7644 52082 7648
rect 52018 7588 52022 7644
rect 52022 7588 52078 7644
rect 52078 7588 52082 7644
rect 52018 7584 52082 7588
rect 52098 7644 52162 7648
rect 52098 7588 52102 7644
rect 52102 7588 52158 7644
rect 52158 7588 52162 7644
rect 52098 7584 52162 7588
rect 21314 7100 21378 7104
rect 21314 7044 21318 7100
rect 21318 7044 21374 7100
rect 21374 7044 21378 7100
rect 21314 7040 21378 7044
rect 21394 7100 21458 7104
rect 21394 7044 21398 7100
rect 21398 7044 21454 7100
rect 21454 7044 21458 7100
rect 21394 7040 21458 7044
rect 21474 7100 21538 7104
rect 21474 7044 21478 7100
rect 21478 7044 21534 7100
rect 21534 7044 21538 7100
rect 21474 7040 21538 7044
rect 21554 7100 21618 7104
rect 21554 7044 21558 7100
rect 21558 7044 21614 7100
rect 21614 7044 21618 7100
rect 21554 7040 21618 7044
rect 41677 7100 41741 7104
rect 41677 7044 41681 7100
rect 41681 7044 41737 7100
rect 41737 7044 41741 7100
rect 41677 7040 41741 7044
rect 41757 7100 41821 7104
rect 41757 7044 41761 7100
rect 41761 7044 41817 7100
rect 41817 7044 41821 7100
rect 41757 7040 41821 7044
rect 41837 7100 41901 7104
rect 41837 7044 41841 7100
rect 41841 7044 41897 7100
rect 41897 7044 41901 7100
rect 41837 7040 41901 7044
rect 41917 7100 41981 7104
rect 41917 7044 41921 7100
rect 41921 7044 41977 7100
rect 41977 7044 41981 7100
rect 41917 7040 41981 7044
rect 11133 6556 11197 6560
rect 11133 6500 11137 6556
rect 11137 6500 11193 6556
rect 11193 6500 11197 6556
rect 11133 6496 11197 6500
rect 11213 6556 11277 6560
rect 11213 6500 11217 6556
rect 11217 6500 11273 6556
rect 11273 6500 11277 6556
rect 11213 6496 11277 6500
rect 11293 6556 11357 6560
rect 11293 6500 11297 6556
rect 11297 6500 11353 6556
rect 11353 6500 11357 6556
rect 11293 6496 11357 6500
rect 11373 6556 11437 6560
rect 11373 6500 11377 6556
rect 11377 6500 11433 6556
rect 11433 6500 11437 6556
rect 11373 6496 11437 6500
rect 31496 6556 31560 6560
rect 31496 6500 31500 6556
rect 31500 6500 31556 6556
rect 31556 6500 31560 6556
rect 31496 6496 31560 6500
rect 31576 6556 31640 6560
rect 31576 6500 31580 6556
rect 31580 6500 31636 6556
rect 31636 6500 31640 6556
rect 31576 6496 31640 6500
rect 31656 6556 31720 6560
rect 31656 6500 31660 6556
rect 31660 6500 31716 6556
rect 31716 6500 31720 6556
rect 31656 6496 31720 6500
rect 31736 6556 31800 6560
rect 31736 6500 31740 6556
rect 31740 6500 31796 6556
rect 31796 6500 31800 6556
rect 31736 6496 31800 6500
rect 51858 6556 51922 6560
rect 51858 6500 51862 6556
rect 51862 6500 51918 6556
rect 51918 6500 51922 6556
rect 51858 6496 51922 6500
rect 51938 6556 52002 6560
rect 51938 6500 51942 6556
rect 51942 6500 51998 6556
rect 51998 6500 52002 6556
rect 51938 6496 52002 6500
rect 52018 6556 52082 6560
rect 52018 6500 52022 6556
rect 52022 6500 52078 6556
rect 52078 6500 52082 6556
rect 52018 6496 52082 6500
rect 52098 6556 52162 6560
rect 52098 6500 52102 6556
rect 52102 6500 52158 6556
rect 52158 6500 52162 6556
rect 52098 6496 52162 6500
rect 21314 6012 21378 6016
rect 21314 5956 21318 6012
rect 21318 5956 21374 6012
rect 21374 5956 21378 6012
rect 21314 5952 21378 5956
rect 21394 6012 21458 6016
rect 21394 5956 21398 6012
rect 21398 5956 21454 6012
rect 21454 5956 21458 6012
rect 21394 5952 21458 5956
rect 21474 6012 21538 6016
rect 21474 5956 21478 6012
rect 21478 5956 21534 6012
rect 21534 5956 21538 6012
rect 21474 5952 21538 5956
rect 21554 6012 21618 6016
rect 21554 5956 21558 6012
rect 21558 5956 21614 6012
rect 21614 5956 21618 6012
rect 21554 5952 21618 5956
rect 41677 6012 41741 6016
rect 41677 5956 41681 6012
rect 41681 5956 41737 6012
rect 41737 5956 41741 6012
rect 41677 5952 41741 5956
rect 41757 6012 41821 6016
rect 41757 5956 41761 6012
rect 41761 5956 41817 6012
rect 41817 5956 41821 6012
rect 41757 5952 41821 5956
rect 41837 6012 41901 6016
rect 41837 5956 41841 6012
rect 41841 5956 41897 6012
rect 41897 5956 41901 6012
rect 41837 5952 41901 5956
rect 41917 6012 41981 6016
rect 41917 5956 41921 6012
rect 41921 5956 41977 6012
rect 41977 5956 41981 6012
rect 41917 5952 41981 5956
rect 37228 5476 37292 5540
rect 11133 5468 11197 5472
rect 11133 5412 11137 5468
rect 11137 5412 11193 5468
rect 11193 5412 11197 5468
rect 11133 5408 11197 5412
rect 11213 5468 11277 5472
rect 11213 5412 11217 5468
rect 11217 5412 11273 5468
rect 11273 5412 11277 5468
rect 11213 5408 11277 5412
rect 11293 5468 11357 5472
rect 11293 5412 11297 5468
rect 11297 5412 11353 5468
rect 11353 5412 11357 5468
rect 11293 5408 11357 5412
rect 11373 5468 11437 5472
rect 11373 5412 11377 5468
rect 11377 5412 11433 5468
rect 11433 5412 11437 5468
rect 11373 5408 11437 5412
rect 31496 5468 31560 5472
rect 31496 5412 31500 5468
rect 31500 5412 31556 5468
rect 31556 5412 31560 5468
rect 31496 5408 31560 5412
rect 31576 5468 31640 5472
rect 31576 5412 31580 5468
rect 31580 5412 31636 5468
rect 31636 5412 31640 5468
rect 31576 5408 31640 5412
rect 31656 5468 31720 5472
rect 31656 5412 31660 5468
rect 31660 5412 31716 5468
rect 31716 5412 31720 5468
rect 31656 5408 31720 5412
rect 31736 5468 31800 5472
rect 31736 5412 31740 5468
rect 31740 5412 31796 5468
rect 31796 5412 31800 5468
rect 31736 5408 31800 5412
rect 51858 5468 51922 5472
rect 51858 5412 51862 5468
rect 51862 5412 51918 5468
rect 51918 5412 51922 5468
rect 51858 5408 51922 5412
rect 51938 5468 52002 5472
rect 51938 5412 51942 5468
rect 51942 5412 51998 5468
rect 51998 5412 52002 5468
rect 51938 5408 52002 5412
rect 52018 5468 52082 5472
rect 52018 5412 52022 5468
rect 52022 5412 52078 5468
rect 52078 5412 52082 5468
rect 52018 5408 52082 5412
rect 52098 5468 52162 5472
rect 52098 5412 52102 5468
rect 52102 5412 52158 5468
rect 52158 5412 52162 5468
rect 52098 5408 52162 5412
rect 37228 5068 37292 5132
rect 21314 4924 21378 4928
rect 21314 4868 21318 4924
rect 21318 4868 21374 4924
rect 21374 4868 21378 4924
rect 21314 4864 21378 4868
rect 21394 4924 21458 4928
rect 21394 4868 21398 4924
rect 21398 4868 21454 4924
rect 21454 4868 21458 4924
rect 21394 4864 21458 4868
rect 21474 4924 21538 4928
rect 21474 4868 21478 4924
rect 21478 4868 21534 4924
rect 21534 4868 21538 4924
rect 21474 4864 21538 4868
rect 21554 4924 21618 4928
rect 21554 4868 21558 4924
rect 21558 4868 21614 4924
rect 21614 4868 21618 4924
rect 21554 4864 21618 4868
rect 41677 4924 41741 4928
rect 41677 4868 41681 4924
rect 41681 4868 41737 4924
rect 41737 4868 41741 4924
rect 41677 4864 41741 4868
rect 41757 4924 41821 4928
rect 41757 4868 41761 4924
rect 41761 4868 41817 4924
rect 41817 4868 41821 4924
rect 41757 4864 41821 4868
rect 41837 4924 41901 4928
rect 41837 4868 41841 4924
rect 41841 4868 41897 4924
rect 41897 4868 41901 4924
rect 41837 4864 41901 4868
rect 41917 4924 41981 4928
rect 41917 4868 41921 4924
rect 41921 4868 41977 4924
rect 41977 4868 41981 4924
rect 41917 4864 41981 4868
rect 11133 4380 11197 4384
rect 11133 4324 11137 4380
rect 11137 4324 11193 4380
rect 11193 4324 11197 4380
rect 11133 4320 11197 4324
rect 11213 4380 11277 4384
rect 11213 4324 11217 4380
rect 11217 4324 11273 4380
rect 11273 4324 11277 4380
rect 11213 4320 11277 4324
rect 11293 4380 11357 4384
rect 11293 4324 11297 4380
rect 11297 4324 11353 4380
rect 11353 4324 11357 4380
rect 11293 4320 11357 4324
rect 11373 4380 11437 4384
rect 11373 4324 11377 4380
rect 11377 4324 11433 4380
rect 11433 4324 11437 4380
rect 11373 4320 11437 4324
rect 31496 4380 31560 4384
rect 31496 4324 31500 4380
rect 31500 4324 31556 4380
rect 31556 4324 31560 4380
rect 31496 4320 31560 4324
rect 31576 4380 31640 4384
rect 31576 4324 31580 4380
rect 31580 4324 31636 4380
rect 31636 4324 31640 4380
rect 31576 4320 31640 4324
rect 31656 4380 31720 4384
rect 31656 4324 31660 4380
rect 31660 4324 31716 4380
rect 31716 4324 31720 4380
rect 31656 4320 31720 4324
rect 31736 4380 31800 4384
rect 31736 4324 31740 4380
rect 31740 4324 31796 4380
rect 31796 4324 31800 4380
rect 31736 4320 31800 4324
rect 51858 4380 51922 4384
rect 51858 4324 51862 4380
rect 51862 4324 51918 4380
rect 51918 4324 51922 4380
rect 51858 4320 51922 4324
rect 51938 4380 52002 4384
rect 51938 4324 51942 4380
rect 51942 4324 51998 4380
rect 51998 4324 52002 4380
rect 51938 4320 52002 4324
rect 52018 4380 52082 4384
rect 52018 4324 52022 4380
rect 52022 4324 52078 4380
rect 52078 4324 52082 4380
rect 52018 4320 52082 4324
rect 52098 4380 52162 4384
rect 52098 4324 52102 4380
rect 52102 4324 52158 4380
rect 52158 4324 52162 4380
rect 52098 4320 52162 4324
rect 21314 3836 21378 3840
rect 21314 3780 21318 3836
rect 21318 3780 21374 3836
rect 21374 3780 21378 3836
rect 21314 3776 21378 3780
rect 21394 3836 21458 3840
rect 21394 3780 21398 3836
rect 21398 3780 21454 3836
rect 21454 3780 21458 3836
rect 21394 3776 21458 3780
rect 21474 3836 21538 3840
rect 21474 3780 21478 3836
rect 21478 3780 21534 3836
rect 21534 3780 21538 3836
rect 21474 3776 21538 3780
rect 21554 3836 21618 3840
rect 21554 3780 21558 3836
rect 21558 3780 21614 3836
rect 21614 3780 21618 3836
rect 21554 3776 21618 3780
rect 41677 3836 41741 3840
rect 41677 3780 41681 3836
rect 41681 3780 41737 3836
rect 41737 3780 41741 3836
rect 41677 3776 41741 3780
rect 41757 3836 41821 3840
rect 41757 3780 41761 3836
rect 41761 3780 41817 3836
rect 41817 3780 41821 3836
rect 41757 3776 41821 3780
rect 41837 3836 41901 3840
rect 41837 3780 41841 3836
rect 41841 3780 41897 3836
rect 41897 3780 41901 3836
rect 41837 3776 41901 3780
rect 41917 3836 41981 3840
rect 41917 3780 41921 3836
rect 41921 3780 41977 3836
rect 41977 3780 41981 3836
rect 41917 3776 41981 3780
rect 11133 3292 11197 3296
rect 11133 3236 11137 3292
rect 11137 3236 11193 3292
rect 11193 3236 11197 3292
rect 11133 3232 11197 3236
rect 11213 3292 11277 3296
rect 11213 3236 11217 3292
rect 11217 3236 11273 3292
rect 11273 3236 11277 3292
rect 11213 3232 11277 3236
rect 11293 3292 11357 3296
rect 11293 3236 11297 3292
rect 11297 3236 11353 3292
rect 11353 3236 11357 3292
rect 11293 3232 11357 3236
rect 11373 3292 11437 3296
rect 11373 3236 11377 3292
rect 11377 3236 11433 3292
rect 11433 3236 11437 3292
rect 11373 3232 11437 3236
rect 31496 3292 31560 3296
rect 31496 3236 31500 3292
rect 31500 3236 31556 3292
rect 31556 3236 31560 3292
rect 31496 3232 31560 3236
rect 31576 3292 31640 3296
rect 31576 3236 31580 3292
rect 31580 3236 31636 3292
rect 31636 3236 31640 3292
rect 31576 3232 31640 3236
rect 31656 3292 31720 3296
rect 31656 3236 31660 3292
rect 31660 3236 31716 3292
rect 31716 3236 31720 3292
rect 31656 3232 31720 3236
rect 31736 3292 31800 3296
rect 31736 3236 31740 3292
rect 31740 3236 31796 3292
rect 31796 3236 31800 3292
rect 31736 3232 31800 3236
rect 51858 3292 51922 3296
rect 51858 3236 51862 3292
rect 51862 3236 51918 3292
rect 51918 3236 51922 3292
rect 51858 3232 51922 3236
rect 51938 3292 52002 3296
rect 51938 3236 51942 3292
rect 51942 3236 51998 3292
rect 51998 3236 52002 3292
rect 51938 3232 52002 3236
rect 52018 3292 52082 3296
rect 52018 3236 52022 3292
rect 52022 3236 52078 3292
rect 52078 3236 52082 3292
rect 52018 3232 52082 3236
rect 52098 3292 52162 3296
rect 52098 3236 52102 3292
rect 52102 3236 52158 3292
rect 52158 3236 52162 3292
rect 52098 3232 52162 3236
rect 21314 2748 21378 2752
rect 21314 2692 21318 2748
rect 21318 2692 21374 2748
rect 21374 2692 21378 2748
rect 21314 2688 21378 2692
rect 21394 2748 21458 2752
rect 21394 2692 21398 2748
rect 21398 2692 21454 2748
rect 21454 2692 21458 2748
rect 21394 2688 21458 2692
rect 21474 2748 21538 2752
rect 21474 2692 21478 2748
rect 21478 2692 21534 2748
rect 21534 2692 21538 2748
rect 21474 2688 21538 2692
rect 21554 2748 21618 2752
rect 21554 2692 21558 2748
rect 21558 2692 21614 2748
rect 21614 2692 21618 2748
rect 21554 2688 21618 2692
rect 41677 2748 41741 2752
rect 41677 2692 41681 2748
rect 41681 2692 41737 2748
rect 41737 2692 41741 2748
rect 41677 2688 41741 2692
rect 41757 2748 41821 2752
rect 41757 2692 41761 2748
rect 41761 2692 41817 2748
rect 41817 2692 41821 2748
rect 41757 2688 41821 2692
rect 41837 2748 41901 2752
rect 41837 2692 41841 2748
rect 41841 2692 41897 2748
rect 41897 2692 41901 2748
rect 41837 2688 41901 2692
rect 41917 2748 41981 2752
rect 41917 2692 41921 2748
rect 41921 2692 41977 2748
rect 41977 2692 41981 2748
rect 41917 2688 41981 2692
rect 11133 2204 11197 2208
rect 11133 2148 11137 2204
rect 11137 2148 11193 2204
rect 11193 2148 11197 2204
rect 11133 2144 11197 2148
rect 11213 2204 11277 2208
rect 11213 2148 11217 2204
rect 11217 2148 11273 2204
rect 11273 2148 11277 2204
rect 11213 2144 11277 2148
rect 11293 2204 11357 2208
rect 11293 2148 11297 2204
rect 11297 2148 11353 2204
rect 11353 2148 11357 2204
rect 11293 2144 11357 2148
rect 11373 2204 11437 2208
rect 11373 2148 11377 2204
rect 11377 2148 11433 2204
rect 11433 2148 11437 2204
rect 11373 2144 11437 2148
rect 31496 2204 31560 2208
rect 31496 2148 31500 2204
rect 31500 2148 31556 2204
rect 31556 2148 31560 2204
rect 31496 2144 31560 2148
rect 31576 2204 31640 2208
rect 31576 2148 31580 2204
rect 31580 2148 31636 2204
rect 31636 2148 31640 2204
rect 31576 2144 31640 2148
rect 31656 2204 31720 2208
rect 31656 2148 31660 2204
rect 31660 2148 31716 2204
rect 31716 2148 31720 2204
rect 31656 2144 31720 2148
rect 31736 2204 31800 2208
rect 31736 2148 31740 2204
rect 31740 2148 31796 2204
rect 31796 2148 31800 2204
rect 31736 2144 31800 2148
rect 51858 2204 51922 2208
rect 51858 2148 51862 2204
rect 51862 2148 51918 2204
rect 51918 2148 51922 2204
rect 51858 2144 51922 2148
rect 51938 2204 52002 2208
rect 51938 2148 51942 2204
rect 51942 2148 51998 2204
rect 51998 2148 52002 2204
rect 51938 2144 52002 2148
rect 52018 2204 52082 2208
rect 52018 2148 52022 2204
rect 52022 2148 52078 2204
rect 52078 2148 52082 2204
rect 52018 2144 52082 2148
rect 52098 2204 52162 2208
rect 52098 2148 52102 2204
rect 52102 2148 52158 2204
rect 52158 2148 52162 2204
rect 52098 2144 52162 2148
<< metal4 >>
rect 11125 17440 11445 17456
rect 11125 17376 11133 17440
rect 11197 17376 11213 17440
rect 11277 17376 11293 17440
rect 11357 17376 11373 17440
rect 11437 17376 11445 17440
rect 11125 16352 11445 17376
rect 11125 16288 11133 16352
rect 11197 16288 11213 16352
rect 11277 16288 11293 16352
rect 11357 16288 11373 16352
rect 11437 16288 11445 16352
rect 11125 15264 11445 16288
rect 11125 15200 11133 15264
rect 11197 15200 11213 15264
rect 11277 15200 11293 15264
rect 11357 15200 11373 15264
rect 11437 15200 11445 15264
rect 11125 14176 11445 15200
rect 11125 14112 11133 14176
rect 11197 14112 11213 14176
rect 11277 14112 11293 14176
rect 11357 14112 11373 14176
rect 11437 14112 11445 14176
rect 11125 13088 11445 14112
rect 11125 13024 11133 13088
rect 11197 13024 11213 13088
rect 11277 13024 11293 13088
rect 11357 13024 11373 13088
rect 11437 13024 11445 13088
rect 11125 12000 11445 13024
rect 11125 11936 11133 12000
rect 11197 11936 11213 12000
rect 11277 11936 11293 12000
rect 11357 11936 11373 12000
rect 11437 11936 11445 12000
rect 11125 10912 11445 11936
rect 11125 10848 11133 10912
rect 11197 10848 11213 10912
rect 11277 10848 11293 10912
rect 11357 10848 11373 10912
rect 11437 10848 11445 10912
rect 11125 9824 11445 10848
rect 11125 9760 11133 9824
rect 11197 9760 11213 9824
rect 11277 9760 11293 9824
rect 11357 9760 11373 9824
rect 11437 9760 11445 9824
rect 11125 8736 11445 9760
rect 11125 8672 11133 8736
rect 11197 8672 11213 8736
rect 11277 8672 11293 8736
rect 11357 8672 11373 8736
rect 11437 8672 11445 8736
rect 11125 7648 11445 8672
rect 11125 7584 11133 7648
rect 11197 7584 11213 7648
rect 11277 7584 11293 7648
rect 11357 7584 11373 7648
rect 11437 7584 11445 7648
rect 11125 6560 11445 7584
rect 11125 6496 11133 6560
rect 11197 6496 11213 6560
rect 11277 6496 11293 6560
rect 11357 6496 11373 6560
rect 11437 6496 11445 6560
rect 11125 5472 11445 6496
rect 11125 5408 11133 5472
rect 11197 5408 11213 5472
rect 11277 5408 11293 5472
rect 11357 5408 11373 5472
rect 11437 5408 11445 5472
rect 11125 4384 11445 5408
rect 11125 4320 11133 4384
rect 11197 4320 11213 4384
rect 11277 4320 11293 4384
rect 11357 4320 11373 4384
rect 11437 4320 11445 4384
rect 11125 3296 11445 4320
rect 11125 3232 11133 3296
rect 11197 3232 11213 3296
rect 11277 3232 11293 3296
rect 11357 3232 11373 3296
rect 11437 3232 11445 3296
rect 11125 2208 11445 3232
rect 11125 2144 11133 2208
rect 11197 2144 11213 2208
rect 11277 2144 11293 2208
rect 11357 2144 11373 2208
rect 11437 2144 11445 2208
rect 11125 2128 11445 2144
rect 21306 16896 21627 17456
rect 21306 16832 21314 16896
rect 21378 16832 21394 16896
rect 21458 16832 21474 16896
rect 21538 16832 21554 16896
rect 21618 16832 21627 16896
rect 21306 15808 21627 16832
rect 21306 15744 21314 15808
rect 21378 15744 21394 15808
rect 21458 15744 21474 15808
rect 21538 15744 21554 15808
rect 21618 15744 21627 15808
rect 21306 14720 21627 15744
rect 21306 14656 21314 14720
rect 21378 14656 21394 14720
rect 21458 14656 21474 14720
rect 21538 14656 21554 14720
rect 21618 14656 21627 14720
rect 21306 13632 21627 14656
rect 21306 13568 21314 13632
rect 21378 13568 21394 13632
rect 21458 13568 21474 13632
rect 21538 13568 21554 13632
rect 21618 13568 21627 13632
rect 21306 12544 21627 13568
rect 21306 12480 21314 12544
rect 21378 12480 21394 12544
rect 21458 12480 21474 12544
rect 21538 12480 21554 12544
rect 21618 12480 21627 12544
rect 21306 11456 21627 12480
rect 21306 11392 21314 11456
rect 21378 11392 21394 11456
rect 21458 11392 21474 11456
rect 21538 11392 21554 11456
rect 21618 11392 21627 11456
rect 21306 10368 21627 11392
rect 21306 10304 21314 10368
rect 21378 10304 21394 10368
rect 21458 10304 21474 10368
rect 21538 10304 21554 10368
rect 21618 10304 21627 10368
rect 21306 9280 21627 10304
rect 21306 9216 21314 9280
rect 21378 9216 21394 9280
rect 21458 9216 21474 9280
rect 21538 9216 21554 9280
rect 21618 9216 21627 9280
rect 21306 8192 21627 9216
rect 21306 8128 21314 8192
rect 21378 8128 21394 8192
rect 21458 8128 21474 8192
rect 21538 8128 21554 8192
rect 21618 8128 21627 8192
rect 21306 7104 21627 8128
rect 21306 7040 21314 7104
rect 21378 7040 21394 7104
rect 21458 7040 21474 7104
rect 21538 7040 21554 7104
rect 21618 7040 21627 7104
rect 21306 6016 21627 7040
rect 21306 5952 21314 6016
rect 21378 5952 21394 6016
rect 21458 5952 21474 6016
rect 21538 5952 21554 6016
rect 21618 5952 21627 6016
rect 21306 4928 21627 5952
rect 21306 4864 21314 4928
rect 21378 4864 21394 4928
rect 21458 4864 21474 4928
rect 21538 4864 21554 4928
rect 21618 4864 21627 4928
rect 21306 3840 21627 4864
rect 21306 3776 21314 3840
rect 21378 3776 21394 3840
rect 21458 3776 21474 3840
rect 21538 3776 21554 3840
rect 21618 3776 21627 3840
rect 21306 2752 21627 3776
rect 21306 2688 21314 2752
rect 21378 2688 21394 2752
rect 21458 2688 21474 2752
rect 21538 2688 21554 2752
rect 21618 2688 21627 2752
rect 21306 2128 21627 2688
rect 31488 17440 31808 17456
rect 31488 17376 31496 17440
rect 31560 17376 31576 17440
rect 31640 17376 31656 17440
rect 31720 17376 31736 17440
rect 31800 17376 31808 17440
rect 31488 16352 31808 17376
rect 31488 16288 31496 16352
rect 31560 16288 31576 16352
rect 31640 16288 31656 16352
rect 31720 16288 31736 16352
rect 31800 16288 31808 16352
rect 31488 15264 31808 16288
rect 31488 15200 31496 15264
rect 31560 15200 31576 15264
rect 31640 15200 31656 15264
rect 31720 15200 31736 15264
rect 31800 15200 31808 15264
rect 31488 14176 31808 15200
rect 31488 14112 31496 14176
rect 31560 14112 31576 14176
rect 31640 14112 31656 14176
rect 31720 14112 31736 14176
rect 31800 14112 31808 14176
rect 31488 13088 31808 14112
rect 31488 13024 31496 13088
rect 31560 13024 31576 13088
rect 31640 13024 31656 13088
rect 31720 13024 31736 13088
rect 31800 13024 31808 13088
rect 31488 12000 31808 13024
rect 31488 11936 31496 12000
rect 31560 11936 31576 12000
rect 31640 11936 31656 12000
rect 31720 11936 31736 12000
rect 31800 11936 31808 12000
rect 31488 10912 31808 11936
rect 31488 10848 31496 10912
rect 31560 10848 31576 10912
rect 31640 10848 31656 10912
rect 31720 10848 31736 10912
rect 31800 10848 31808 10912
rect 31488 9824 31808 10848
rect 31488 9760 31496 9824
rect 31560 9760 31576 9824
rect 31640 9760 31656 9824
rect 31720 9760 31736 9824
rect 31800 9760 31808 9824
rect 31488 8736 31808 9760
rect 31488 8672 31496 8736
rect 31560 8672 31576 8736
rect 31640 8672 31656 8736
rect 31720 8672 31736 8736
rect 31800 8672 31808 8736
rect 31488 7648 31808 8672
rect 31488 7584 31496 7648
rect 31560 7584 31576 7648
rect 31640 7584 31656 7648
rect 31720 7584 31736 7648
rect 31800 7584 31808 7648
rect 31488 6560 31808 7584
rect 31488 6496 31496 6560
rect 31560 6496 31576 6560
rect 31640 6496 31656 6560
rect 31720 6496 31736 6560
rect 31800 6496 31808 6560
rect 31488 5472 31808 6496
rect 41669 16896 41989 17456
rect 41669 16832 41677 16896
rect 41741 16832 41757 16896
rect 41821 16832 41837 16896
rect 41901 16832 41917 16896
rect 41981 16832 41989 16896
rect 41669 15808 41989 16832
rect 41669 15744 41677 15808
rect 41741 15744 41757 15808
rect 41821 15744 41837 15808
rect 41901 15744 41917 15808
rect 41981 15744 41989 15808
rect 41669 14720 41989 15744
rect 41669 14656 41677 14720
rect 41741 14656 41757 14720
rect 41821 14656 41837 14720
rect 41901 14656 41917 14720
rect 41981 14656 41989 14720
rect 41669 13632 41989 14656
rect 41669 13568 41677 13632
rect 41741 13568 41757 13632
rect 41821 13568 41837 13632
rect 41901 13568 41917 13632
rect 41981 13568 41989 13632
rect 41669 12544 41989 13568
rect 41669 12480 41677 12544
rect 41741 12480 41757 12544
rect 41821 12480 41837 12544
rect 41901 12480 41917 12544
rect 41981 12480 41989 12544
rect 41669 11456 41989 12480
rect 41669 11392 41677 11456
rect 41741 11392 41757 11456
rect 41821 11392 41837 11456
rect 41901 11392 41917 11456
rect 41981 11392 41989 11456
rect 41669 10368 41989 11392
rect 41669 10304 41677 10368
rect 41741 10304 41757 10368
rect 41821 10304 41837 10368
rect 41901 10304 41917 10368
rect 41981 10304 41989 10368
rect 41669 9280 41989 10304
rect 41669 9216 41677 9280
rect 41741 9216 41757 9280
rect 41821 9216 41837 9280
rect 41901 9216 41917 9280
rect 41981 9216 41989 9280
rect 41669 8192 41989 9216
rect 41669 8128 41677 8192
rect 41741 8128 41757 8192
rect 41821 8128 41837 8192
rect 41901 8128 41917 8192
rect 41981 8128 41989 8192
rect 41669 7104 41989 8128
rect 41669 7040 41677 7104
rect 41741 7040 41757 7104
rect 41821 7040 41837 7104
rect 41901 7040 41917 7104
rect 41981 7040 41989 7104
rect 41669 6016 41989 7040
rect 41669 5952 41677 6016
rect 41741 5952 41757 6016
rect 41821 5952 41837 6016
rect 41901 5952 41917 6016
rect 41981 5952 41989 6016
rect 37227 5540 37293 5541
rect 37227 5476 37228 5540
rect 37292 5476 37293 5540
rect 37227 5475 37293 5476
rect 31488 5408 31496 5472
rect 31560 5408 31576 5472
rect 31640 5408 31656 5472
rect 31720 5408 31736 5472
rect 31800 5408 31808 5472
rect 31488 4384 31808 5408
rect 37230 5133 37290 5475
rect 37227 5132 37293 5133
rect 37227 5068 37228 5132
rect 37292 5068 37293 5132
rect 37227 5067 37293 5068
rect 31488 4320 31496 4384
rect 31560 4320 31576 4384
rect 31640 4320 31656 4384
rect 31720 4320 31736 4384
rect 31800 4320 31808 4384
rect 31488 3296 31808 4320
rect 31488 3232 31496 3296
rect 31560 3232 31576 3296
rect 31640 3232 31656 3296
rect 31720 3232 31736 3296
rect 31800 3232 31808 3296
rect 31488 2208 31808 3232
rect 31488 2144 31496 2208
rect 31560 2144 31576 2208
rect 31640 2144 31656 2208
rect 31720 2144 31736 2208
rect 31800 2144 31808 2208
rect 31488 2128 31808 2144
rect 41669 4928 41989 5952
rect 41669 4864 41677 4928
rect 41741 4864 41757 4928
rect 41821 4864 41837 4928
rect 41901 4864 41917 4928
rect 41981 4864 41989 4928
rect 41669 3840 41989 4864
rect 41669 3776 41677 3840
rect 41741 3776 41757 3840
rect 41821 3776 41837 3840
rect 41901 3776 41917 3840
rect 41981 3776 41989 3840
rect 41669 2752 41989 3776
rect 41669 2688 41677 2752
rect 41741 2688 41757 2752
rect 41821 2688 41837 2752
rect 41901 2688 41917 2752
rect 41981 2688 41989 2752
rect 41669 2128 41989 2688
rect 51850 17440 52170 17456
rect 51850 17376 51858 17440
rect 51922 17376 51938 17440
rect 52002 17376 52018 17440
rect 52082 17376 52098 17440
rect 52162 17376 52170 17440
rect 51850 16352 52170 17376
rect 51850 16288 51858 16352
rect 51922 16288 51938 16352
rect 52002 16288 52018 16352
rect 52082 16288 52098 16352
rect 52162 16288 52170 16352
rect 51850 15264 52170 16288
rect 51850 15200 51858 15264
rect 51922 15200 51938 15264
rect 52002 15200 52018 15264
rect 52082 15200 52098 15264
rect 52162 15200 52170 15264
rect 51850 14176 52170 15200
rect 51850 14112 51858 14176
rect 51922 14112 51938 14176
rect 52002 14112 52018 14176
rect 52082 14112 52098 14176
rect 52162 14112 52170 14176
rect 51850 13088 52170 14112
rect 51850 13024 51858 13088
rect 51922 13024 51938 13088
rect 52002 13024 52018 13088
rect 52082 13024 52098 13088
rect 52162 13024 52170 13088
rect 51850 12000 52170 13024
rect 51850 11936 51858 12000
rect 51922 11936 51938 12000
rect 52002 11936 52018 12000
rect 52082 11936 52098 12000
rect 52162 11936 52170 12000
rect 51850 10912 52170 11936
rect 51850 10848 51858 10912
rect 51922 10848 51938 10912
rect 52002 10848 52018 10912
rect 52082 10848 52098 10912
rect 52162 10848 52170 10912
rect 51850 9824 52170 10848
rect 51850 9760 51858 9824
rect 51922 9760 51938 9824
rect 52002 9760 52018 9824
rect 52082 9760 52098 9824
rect 52162 9760 52170 9824
rect 51850 8736 52170 9760
rect 51850 8672 51858 8736
rect 51922 8672 51938 8736
rect 52002 8672 52018 8736
rect 52082 8672 52098 8736
rect 52162 8672 52170 8736
rect 51850 7648 52170 8672
rect 51850 7584 51858 7648
rect 51922 7584 51938 7648
rect 52002 7584 52018 7648
rect 52082 7584 52098 7648
rect 52162 7584 52170 7648
rect 51850 6560 52170 7584
rect 51850 6496 51858 6560
rect 51922 6496 51938 6560
rect 52002 6496 52018 6560
rect 52082 6496 52098 6560
rect 52162 6496 52170 6560
rect 51850 5472 52170 6496
rect 51850 5408 51858 5472
rect 51922 5408 51938 5472
rect 52002 5408 52018 5472
rect 52082 5408 52098 5472
rect 52162 5408 52170 5472
rect 51850 4384 52170 5408
rect 51850 4320 51858 4384
rect 51922 4320 51938 4384
rect 52002 4320 52018 4384
rect 52082 4320 52098 4384
rect 52162 4320 52170 4384
rect 51850 3296 52170 4320
rect 51850 3232 51858 3296
rect 51922 3232 51938 3296
rect 52002 3232 52018 3296
rect 52082 3232 52098 3296
rect 52162 3232 52170 3296
rect 51850 2208 52170 3232
rect 51850 2144 51858 2208
rect 51922 2144 51938 2208
rect 52002 2144 52018 2208
rect 52082 2144 52098 2208
rect 52162 2144 52170 2208
rect 51850 2128 52170 2144
use sky130_fd_sc_hd__decap_12  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1607721120
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 2116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 1380 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1607721120
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1607721120
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0624_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1607721120
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1607721120
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23
timestamp 1607721120
transform 1 0 3220 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1310_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 4324 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _0942_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 4692 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_1_53
timestamp 1607721120
transform 1 0 5980 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54
timestamp 1607721120
transform 1 0 6072 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1607721120
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1607721120
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1309_
timestamp 1607721120
transform 1 0 6900 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__a21boi_4  _0937_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 6808 0 1 2720
box -38 -48 1418 592
use sky130_fd_sc_hd__decap_12  FILLER_1_89
timestamp 1607721120
transform 1 0 9292 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_77
timestamp 1607721120
transform 1 0 8188 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_90
timestamp 1607721120
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82
timestamp 1607721120
transform 1 0 8648 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1607721120
transform 1 0 11500 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_101
timestamp 1607721120
transform 1 0 10396 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1607721120
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1607721120
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1607721120
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1607721120
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1607721120
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1607721120
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1313_
timestamp 1607721120
transform 1 0 12604 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _0917_
timestamp 1607721120
transform 1 0 12696 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_1_152
timestamp 1607721120
transform 1 0 15088 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_140
timestamp 1607721120
transform 1 0 13984 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp 1607721120
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 1607721120
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_144
timestamp 1607721120
transform 1 0 14352 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1607721120
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1314_
timestamp 1607721120
transform 1 0 15732 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0915_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 14720 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_175
timestamp 1607721120
transform 1 0 17204 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_160
timestamp 1607721120
transform 1 0 15824 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_178
timestamp 1607721120
transform 1 0 17480 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0903_
timestamp 1607721120
transform 1 0 15916 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_1_198
timestamp 1607721120
transform 1 0 19320 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1607721120
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1607721120
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1315_
timestamp 1607721120
transform 1 0 18308 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _0912_
timestamp 1607721120
transform 1 0 18032 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_1_218
timestamp 1607721120
transform 1 0 21160 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_227
timestamp 1607721120
transform 1 0 21988 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_214
timestamp 1607721120
transform 1 0 20792 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_206
timestamp 1607721120
transform 1 0 20056 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1607721120
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0900_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _0894_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 20056 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_236
timestamp 1607721120
transform 1 0 22816 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_230 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 22264 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_235
timestamp 1607721120
transform 1 0 22724 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0828_
timestamp 1607721120
transform 1 0 22448 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0827_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 22908 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_245
timestamp 1607721120
transform 1 0 23644 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_240
timestamp 1607721120
transform 1 0 23184 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1607721120
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1607721120
transform 1 0 24012 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1607721120
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_274
timestamp 1607721120
transform 1 0 26312 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_253
timestamp 1607721120
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_271
timestamp 1607721120
transform 1 0 26036 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1323_
timestamp 1607721120
transform 1 0 24288 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1319_
timestamp 1607721120
transform 1 0 24564 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_286
timestamp 1607721120
transform 1 0 27416 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_295
timestamp 1607721120
transform 1 0 28244 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1607721120
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__a21boi_4  _0831_
timestamp 1607721120
transform 1 0 26864 0 -1 2720
box -38 -48 1418 592
use sky130_fd_sc_hd__and3_4  _0816_
timestamp 1607721120
transform 1 0 27600 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_312
timestamp 1607721120
transform 1 0 29808 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_306
timestamp 1607721120
transform 1 0 29256 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_297
timestamp 1607721120
transform 1 0 28428 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_311
timestamp 1607721120
transform 1 0 29716 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_307
timestamp 1607721120
transform 1 0 29348 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1607721120
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1607721120
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1283_
timestamp 1607721120
transform 1 0 29992 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 29900 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_325
timestamp 1607721120
transform 1 0 31004 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_333
timestamp 1607721120
transform 1 0 31740 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1607721120
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1099_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 31740 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _0642_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 32568 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_1_358
timestamp 1607721120
transform 1 0 34040 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_347
timestamp 1607721120
transform 1 0 33028 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_364
timestamp 1607721120
transform 1 0 34592 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_349
timestamp 1607721120
transform 1 0 33212 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0822_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 33948 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1607721120
transform 1 0 33764 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_385
timestamp 1607721120
transform 1 0 36524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_375
timestamp 1607721120
transform 1 0 35604 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_367
timestamp 1607721120
transform 1 0 34868 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_386
timestamp 1607721120
transform 1 0 36616 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1607721120
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1607721120
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0649_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 35696 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_4  _0641_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 35420 0 -1 2720
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_1_397
timestamp 1607721120
transform 1 0 37628 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_404
timestamp 1607721120
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_402
timestamp 1607721120
transform 1 0 38088 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_398 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 37720 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1607721120
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1324_
timestamp 1607721120
transform 1 0 37904 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1281_
timestamp 1607721120
transform 1 0 38548 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_1_419
timestamp 1607721120
transform 1 0 39652 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_426
timestamp 1607721120
transform 1 0 40296 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1607721120
transform 1 0 40388 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0625_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 40480 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_1_448
timestamp 1607721120
transform 1 0 42320 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_437
timestamp 1607721120
transform 1 0 41308 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_455
timestamp 1607721120
transform 1 0 42964 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_444
timestamp 1607721120
transform 1 0 41952 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1607721120
transform 1 0 41032 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1101_
timestamp 1607721120
transform 1 0 42044 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1607721120
transform 1 0 42688 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0623_
timestamp 1607721120
transform 1 0 41124 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_472
timestamp 1607721120
transform 1 0 44528 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_460
timestamp 1607721120
transform 1 0 43424 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_470
timestamp 1607721120
transform 1 0 44344 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_466
timestamp 1607721120
transform 1 0 43976 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_463
timestamp 1607721120
transform 1 0 43700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1607721120
transform 1 0 43884 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0628_
timestamp 1607721120
transform 1 0 44620 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0627_
timestamp 1607721120
transform 1 0 44436 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_1_480
timestamp 1607721120
transform 1 0 45264 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_497
timestamp 1607721120
transform 1 0 46828 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_492
timestamp 1607721120
transform 1 0 46368 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_480
timestamp 1607721120
transform 1 0 45264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1607721120
transform 1 0 46000 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1607721120
transform 1 0 46736 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__nor4_4  _0637_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 46092 0 1 2720
box -38 -48 1602 592
use sky130_fd_sc_hd__or4_4  _0626_
timestamp 1607721120
transform 1 0 46920 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_1_523
timestamp 1607721120
transform 1 0 49220 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_506
timestamp 1607721120
transform 1 0 47656 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_519
timestamp 1607721120
transform 1 0 48852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_507
timestamp 1607721120
transform 1 0 47748 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0653_
timestamp 1607721120
transform 1 0 48484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _0652_
timestamp 1607721120
transform 1 0 48392 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_547
timestamp 1607721120
transform 1 0 51428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_535
timestamp 1607721120
transform 1 0 50324 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_540
timestamp 1607721120
transform 1 0 50784 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_528
timestamp 1607721120
transform 1 0 49680 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1607721120
transform 1 0 49588 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0687_
timestamp 1607721120
transform 1 0 49956 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_560
timestamp 1607721120
transform 1 0 52624 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_550
timestamp 1607721120
transform 1 0 51704 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_559
timestamp 1607721120
transform 1 0 52532 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_552
timestamp 1607721120
transform 1 0 51888 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1607721120
transform 1 0 51612 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1607721120
transform 1 0 52440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1093_
timestamp 1607721120
transform 1 0 53360 0 1 2720
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _0680_
timestamp 1607721120
transform 1 0 52256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_582
timestamp 1607721120
transform 1 0 54648 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_590
timestamp 1607721120
transform 1 0 55384 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_581
timestamp 1607721120
transform 1 0 54556 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_571
timestamp 1607721120
transform 1 0 53636 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1607721120
transform 1 0 55292 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1081_
timestamp 1607721120
transform 1 0 55384 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0630_
timestamp 1607721120
transform 1 0 53728 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_1_611
timestamp 1607721120
transform 1 0 57316 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_609
timestamp 1607721120
transform 1 0 57132 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_597
timestamp 1607721120
transform 1 0 56028 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_612
timestamp 1607721120
transform 1 0 57408 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_602
timestamp 1607721120
transform 1 0 56488 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1607721120
transform 1 0 57224 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0631_
timestamp 1607721120
transform 1 0 56764 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_1_631
timestamp 1607721120
transform 1 0 59156 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_619
timestamp 1607721120
transform 1 0 58052 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_630
timestamp 1607721120
transform 1 0 59064 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1607721120
transform 1 0 58144 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0636_
timestamp 1607721120
transform 1 0 58328 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0635_
timestamp 1607721120
transform 1 0 59892 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0632_
timestamp 1607721120
transform 1 0 58236 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1607721120
transform 1 0 59800 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_658
timestamp 1607721120
transform 1 0 61640 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_646
timestamp 1607721120
transform 1 0 60536 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_660
timestamp 1607721120
transform 1 0 61824 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_652
timestamp 1607721120
transform 1 0 61088 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_649
timestamp 1607721120
transform 1 0 60812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_641
timestamp 1607721120
transform 1 0 60076 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1607721120
transform 1 0 60996 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1607721120
transform -1 0 62192 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1607721120
transform -1 0 62192 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1607721120
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1607721120
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1607721120
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_43
timestamp 1607721120
transform 1 0 5060 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1607721120
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1607721120
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1607721120
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0941_
timestamp 1607721120
transform 1 0 4416 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_2_65
timestamp 1607721120
transform 1 0 7084 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0938_
timestamp 1607721120
transform 1 0 5796 0 -1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1607721120
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_82
timestamp 1607721120
transform 1 0 8648 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _0936_
timestamp 1607721120
transform 1 0 7820 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1607721120
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1607721120
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1607721120
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_137
timestamp 1607721120
transform 1 0 13708 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_122
timestamp 1607721120
transform 1 0 12328 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_117
timestamp 1607721120
transform 1 0 11868 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0913_
timestamp 1607721120
transform 1 0 13064 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0789_
timestamp 1607721120
transform 1 0 11960 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_154
timestamp 1607721120
transform 1 0 15272 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1607721120
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1607721120
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_181
timestamp 1607721120
transform 1 0 17756 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_162
timestamp 1607721120
transform 1 0 16008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _0914_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 16284 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1607721120
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _0899_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 18492 0 -1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_2_219
timestamp 1607721120
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1607721120
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0897_
timestamp 1607721120
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_247
timestamp 1607721120
transform 1 0 23828 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_239
timestamp 1607721120
transform 1 0 23092 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_231
timestamp 1607721120
transform 1 0 22356 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0943_
timestamp 1607721120
transform 1 0 23184 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_2_267
timestamp 1607721120
transform 1 0 25668 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _0852_
timestamp 1607721120
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_296
timestamp 1607721120
transform 1 0 28336 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_284
timestamp 1607721120
transform 1 0 27232 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_276
timestamp 1607721120
transform 1 0 26496 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1607721120
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0829_
timestamp 1607721120
transform 1 0 27508 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_319
timestamp 1607721120
transform 1 0 30452 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_308
timestamp 1607721120
transform 1 0 29440 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0832_
timestamp 1607721120
transform 1 0 29624 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_335
timestamp 1607721120
transform 1 0 31924 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_331
timestamp 1607721120
transform 1 0 31556 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1607721120
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1098_
timestamp 1607721120
transform 1 0 32108 0 -1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_2_351
timestamp 1607721120
transform 1 0 33396 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _0840_
timestamp 1607721120
transform 1 0 34132 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_385
timestamp 1607721120
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_368
timestamp 1607721120
transform 1 0 34960 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 35512 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1102_
timestamp 1607721120
transform 1 0 35696 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_410
timestamp 1607721120
transform 1 0 38824 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_402
timestamp 1607721120
transform 1 0 38088 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1607721120
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1321_
timestamp 1607721120
transform 1 0 38916 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0895_
timestamp 1607721120
transform 1 0 37720 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_430
timestamp 1607721120
transform 1 0 40664 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_454
timestamp 1607721120
transform 1 0 42872 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_442
timestamp 1607721120
transform 1 0 41768 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0935_
timestamp 1607721120
transform 1 0 41400 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_471
timestamp 1607721120
transform 1 0 44436 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_459
timestamp 1607721120
transform 1 0 43332 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1607721120
transform 1 0 43240 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0638_
timestamp 1607721120
transform 1 0 45172 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_483
timestamp 1607721120
transform 1 0 45540 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1284_
timestamp 1607721120
transform 1 0 46276 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_2_520
timestamp 1607721120
transform 1 0 48944 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_518
timestamp 1607721120
transform 1 0 48760 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_510
timestamp 1607721120
transform 1 0 48024 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1607721120
transform 1 0 48852 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_546
timestamp 1607721120
transform 1 0 51336 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_534
timestamp 1607721120
transform 1 0 50232 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_526
timestamp 1607721120
transform 1 0 49496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1092_
timestamp 1607721120
transform 1 0 51520 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1084_
timestamp 1607721120
transform 1 0 49588 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_2_555
timestamp 1607721120
transform 1 0 52164 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0634_
timestamp 1607721120
transform 1 0 52900 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_581
timestamp 1607721120
transform 1 0 54556 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_572
timestamp 1607721120
transform 1 0 53728 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1607721120
transform 1 0 54464 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1091_
timestamp 1607721120
transform 1 0 54648 0 -1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_2_611
timestamp 1607721120
transform 1 0 57316 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_596
timestamp 1607721120
transform 1 0 55936 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1090_
timestamp 1607721120
transform 1 0 56672 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_2_633
timestamp 1607721120
transform 1 0 59340 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1089_
timestamp 1607721120
transform 1 0 58052 0 -1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_2_657
timestamp 1607721120
transform 1 0 61548 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_645
timestamp 1607721120
transform 1 0 60444 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1607721120
transform 1 0 60076 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1607721120
transform -1 0 62192 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1607721120
transform 1 0 60168 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp 1607721120
transform 1 0 2484 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1607721120
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1607721120
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1167_
timestamp 1607721120
transform 1 0 2576 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_3_38
timestamp 1607721120
transform 1 0 4600 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_23
timestamp 1607721120
transform 1 0 3220 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1165_
timestamp 1607721120
transform 1 0 3956 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_3_53
timestamp 1607721120
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1607721120
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0940_
timestamp 1607721120
transform 1 0 6808 0 1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _0939_
timestamp 1607721120
transform 1 0 5336 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_3_88
timestamp 1607721120
transform 1 0 9200 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_76
timestamp 1607721120
transform 1 0 8096 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0809_
timestamp 1607721120
transform 1 0 8832 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_112
timestamp 1607721120
transform 1 0 11408 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_100
timestamp 1607721120
transform 1 0 10304 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_137
timestamp 1607721120
transform 1 0 13708 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_129
timestamp 1607721120
transform 1 0 12972 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_123
timestamp 1607721120
transform 1 0 12420 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1607721120
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1607721120
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0916_
timestamp 1607721120
transform 1 0 13064 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_3_155
timestamp 1607721120
transform 1 0 15364 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_145
timestamp 1607721120
transform 1 0 14444 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0883_
timestamp 1607721120
transform 1 0 14720 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_3_175
timestamp 1607721120
transform 1 0 17204 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _0911_
timestamp 1607721120
transform 1 0 16100 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_198
timestamp 1607721120
transform 1 0 19320 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_184
timestamp 1607721120
transform 1 0 18032 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1607721120
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_4  _0908_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 18124 0 1 3808
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_3_227
timestamp 1607721120
transform 1 0 21988 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_215
timestamp 1607721120
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_4  _1187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 20056 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_245
timestamp 1607721120
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_236
timestamp 1607721120
transform 1 0 22816 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_231
timestamp 1607721120
transform 1 0 22356 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1607721120
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0851_
timestamp 1607721120
transform 1 0 22448 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _0850_
timestamp 1607721120
transform 1 0 23736 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_3_273
timestamp 1607721120
transform 1 0 26220 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_253
timestamp 1607721120
transform 1 0 24380 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _0830_
timestamp 1607721120
transform 1 0 25116 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_288
timestamp 1607721120
transform 1 0 27600 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1244_
timestamp 1607721120
transform 1 0 26956 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_3_312
timestamp 1607721120
transform 1 0 29808 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_306
timestamp 1607721120
transform 1 0 29256 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_304
timestamp 1607721120
transform 1 0 29072 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_300
timestamp 1607721120
transform 1 0 28704 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1607721120
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1100_
timestamp 1607721120
transform 1 0 29900 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_322
timestamp 1607721120
transform 1 0 30728 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1320_
timestamp 1607721120
transform 1 0 31464 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_3_365
timestamp 1607721120
transform 1 0 34684 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_361
timestamp 1607721120
transform 1 0 34316 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1607721120
transform 1 0 33212 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_382
timestamp 1607721120
transform 1 0 36248 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_371
timestamp 1607721120
transform 1 0 35236 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1607721120
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0863_
timestamp 1607721120
transform 1 0 34868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1607721120
transform 1 0 35972 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_399
timestamp 1607721120
transform 1 0 37812 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _0846_
timestamp 1607721120
transform 1 0 38548 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _0826_
timestamp 1607721120
transform 1 0 36984 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_428
timestamp 1607721120
transform 1 0 40480 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_419
timestamp 1607721120
transform 1 0 39652 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1607721120
transform 1 0 40388 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1322_
timestamp 1607721120
transform 1 0 40572 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_3_448
timestamp 1607721120
transform 1 0 42320 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_468
timestamp 1607721120
transform 1 0 44160 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_460
timestamp 1607721120
transform 1 0 43424 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1103_
timestamp 1607721120
transform 1 0 43792 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0905_
timestamp 1607721120
transform 1 0 44896 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_489
timestamp 1607721120
transform 1 0 46092 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_480
timestamp 1607721120
transform 1 0 45264 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1607721120
transform 1 0 46000 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1097_
timestamp 1607721120
transform 1 0 46460 0 1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_3_519
timestamp 1607721120
transform 1 0 48852 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_507
timestamp 1607721120
transform 1 0 47748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _1085_
timestamp 1607721120
transform 1 0 49128 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_546
timestamp 1607721120
transform 1 0 51336 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_534
timestamp 1607721120
transform 1 0 50232 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_550
timestamp 1607721120
transform 1 0 51704 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1607721120
transform 1 0 51612 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1285_
timestamp 1607721120
transform 1 0 52256 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_3_575
timestamp 1607721120
transform 1 0 54004 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _1087_
timestamp 1607721120
transform 1 0 55108 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_616
timestamp 1607721120
transform 1 0 57776 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_611
timestamp 1607721120
transform 1 0 57316 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_608
timestamp 1607721120
transform 1 0 57040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_596
timestamp 1607721120
transform 1 0 55936 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1607721120
transform 1 0 57224 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1070_
timestamp 1607721120
transform 1 0 57408 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1286_
timestamp 1607721120
transform 1 0 58512 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_3_655
timestamp 1607721120
transform 1 0 61364 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_643
timestamp 1607721120
transform 1 0 60260 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1607721120
transform -1 0 62192 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_15
timestamp 1607721120
transform 1 0 2484 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1607721120
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1607721120
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1169_
timestamp 1607721120
transform 1 0 2576 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_4_43
timestamp 1607721120
transform 1 0 5060 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_35
timestamp 1607721120
transform 1 0 4324 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_23
timestamp 1607721120
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1607721120
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1188_
timestamp 1607721120
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_58
timestamp 1607721120
transform 1 0 6440 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_4  _0934_
timestamp 1607721120
transform 1 0 7176 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_4  _0933_
timestamp 1607721120
transform 1 0 5336 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1607721120
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_79
timestamp 1607721120
transform 1 0 8372 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_113
timestamp 1607721120
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_105
timestamp 1607721120
transform 1 0 10764 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1607721120
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1607721120
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_124
timestamp 1607721120
transform 1 0 12512 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _0889_
timestamp 1607721120
transform 1 0 13248 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0884_
timestamp 1607721120
transform 1 0 11684 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1607721120
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1607721120
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0885_
timestamp 1607721120
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_163
timestamp 1607721120
transform 1 0 16100 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _0910_
timestamp 1607721120
transform 1 0 16836 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_200
timestamp 1607721120
transform 1 0 19504 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_183
timestamp 1607721120
transform 1 0 17940 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _0919_
timestamp 1607721120
transform 1 0 18676 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_223
timestamp 1607721120
transform 1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1607721120
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1607721120
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1607721120
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _0892_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 21896 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_4_247
timestamp 1607721120
transform 1 0 23828 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_239
timestamp 1607721120
transform 1 0 23092 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_4  _0896_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 24104 0 -1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_4_267
timestamp 1607721120
transform 1 0 25668 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_283
timestamp 1607721120
transform 1 0 27140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1607721120
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0818_
timestamp 1607721120
transform 1 0 28244 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _0815_
timestamp 1607721120
transform 1 0 26496 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_4_304
timestamp 1607721120
transform 1 0 29072 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _0849_
timestamp 1607721120
transform 1 0 30176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_328
timestamp 1607721120
transform 1 0 31280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1607721120
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1282_
timestamp 1607721120
transform 1 0 32108 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_4_356
timestamp 1607721120
transform 1 0 33856 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_374
timestamp 1607721120
transform 1 0 35512 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_368
timestamp 1607721120
transform 1 0 34960 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0825_
timestamp 1607721120
transform 1 0 36248 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0741_
timestamp 1607721120
transform 1 0 35144 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_402
timestamp 1607721120
transform 1 0 38088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_398
timestamp 1607721120
transform 1 0 37720 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_389
timestamp 1607721120
transform 1 0 36892 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1607721120
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1108_
timestamp 1607721120
transform 1 0 38180 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_428
timestamp 1607721120
transform 1 0 40480 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_424
timestamp 1607721120
transform 1 0 40112 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_412
timestamp 1607721120
transform 1 0 39008 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _0843_
timestamp 1607721120
transform 1 0 40572 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_453
timestamp 1607721120
transform 1 0 42780 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_441
timestamp 1607721120
transform 1 0 41676 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_478
timestamp 1607721120
transform 1 0 45080 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_466
timestamp 1607721120
transform 1 0 43976 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_457
timestamp 1607721120
transform 1 0 43148 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1607721120
transform 1 0 43240 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1074_
timestamp 1607721120
transform 1 0 43332 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_4_500
timestamp 1607721120
transform 1 0 47104 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_485
timestamp 1607721120
transform 1 0 45724 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1153_
timestamp 1607721120
transform 1 0 46460 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0869_
timestamp 1607721120
transform 1 0 45356 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_511
timestamp 1607721120
transform 1 0 48116 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1607721120
transform 1 0 48852 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1287_
timestamp 1607721120
transform 1 0 48944 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1079_
timestamp 1607721120
transform 1 0 47840 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_539
timestamp 1607721120
transform 1 0 50692 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _1083_
timestamp 1607721120
transform 1 0 51428 0 -1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_4_561
timestamp 1607721120
transform 1 0 52716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_589
timestamp 1607721120
transform 1 0 55292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_581
timestamp 1607721120
transform 1 0 54556 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_579
timestamp 1607721120
transform 1 0 54372 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_573
timestamp 1607721120
transform 1 0 53820 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1607721120
transform 1 0 54464 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_4  _1086_
timestamp 1607721120
transform 1 0 55568 0 -1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_4_605
timestamp 1607721120
transform 1 0 56764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_633
timestamp 1607721120
transform 1 0 59340 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_617
timestamp 1607721120
transform 1 0 57868 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a21boi_4  _1088_
timestamp 1607721120
transform 1 0 57960 0 -1 4896
box -38 -48 1418 592
use sky130_fd_sc_hd__fill_1  FILLER_4_660
timestamp 1607721120
transform 1 0 61824 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_654
timestamp 1607721120
transform 1 0 61272 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_642
timestamp 1607721120
transform 1 0 60168 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1607721120
transform 1 0 60076 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1607721120
transform -1 0 62192 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp 1607721120
transform 1 0 2484 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1607721120
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1607721120
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1171_
timestamp 1607721120
transform 1 0 2760 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_5_25
timestamp 1607721120
transform 1 0 3404 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1311_
timestamp 1607721120
transform 1 0 4140 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1607721120
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_52
timestamp 1607721120
transform 1 0 5888 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1607721120
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0931_
timestamp 1607721120
transform 1 0 6808 0 1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_5_91
timestamp 1607721120
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_76
timestamp 1607721120
transform 1 0 8096 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0929_
timestamp 1607721120
transform 1 0 8832 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_5_112
timestamp 1607721120
transform 1 0 11408 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0997_
timestamp 1607721120
transform 1 0 10580 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_137
timestamp 1607721120
transform 1 0 13708 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1607721120
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1607721120
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0947_
timestamp 1607721120
transform 1 0 12420 0 1 4896
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_5_155
timestamp 1607721120
transform 1 0 15364 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_145
timestamp 1607721120
transform 1 0 14444 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0924_
timestamp 1607721120
transform 1 0 14720 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_5_175
timestamp 1607721120
transform 1 0 17204 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _0925_
timestamp 1607721120
transform 1 0 16100 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_193
timestamp 1607721120
transform 1 0 18860 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1607721120
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0926_
timestamp 1607721120
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _0922_
timestamp 1607721120
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1607721120
transform 1 0 21804 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_210
timestamp 1607721120
transform 1 0 20424 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0921_
timestamp 1607721120
transform 1 0 21160 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_5_245
timestamp 1607721120
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_243
timestamp 1607721120
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_237
timestamp 1607721120
transform 1 0 22908 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1607721120
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _0893_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 24012 0 1 4896
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_5_271
timestamp 1607721120
transform 1 0 26036 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_288
timestamp 1607721120
transform 1 0 27600 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _1163_
timestamp 1607721120
transform 1 0 26772 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_314
timestamp 1607721120
transform 1 0 29992 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_306
timestamp 1607721120
transform 1 0 29256 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_304
timestamp 1607721120
transform 1 0 29072 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_300
timestamp 1607721120
transform 1 0 28704 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1607721120
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0643_
timestamp 1607721120
transform 1 0 30268 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_342
timestamp 1607721120
transform 1 0 32568 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_321
timestamp 1607721120
transform 1 0 30636 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _0842_
timestamp 1607721120
transform 1 0 31372 0 1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_5_354
timestamp 1607721120
transform 1 0 33672 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0836_
timestamp 1607721120
transform 1 0 33304 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_370
timestamp 1607721120
transform 1 0 35144 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1607721120
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _1057_
timestamp 1607721120
transform 1 0 35880 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1607721120
transform 1 0 34868 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_411
timestamp 1607721120
transform 1 0 38916 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_407
timestamp 1607721120
transform 1 0 38548 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_395
timestamp 1607721120
transform 1 0 37444 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_428
timestamp 1607721120
transform 1 0 40480 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_419
timestamp 1607721120
transform 1 0 39652 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1607721120
transform 1 0 40388 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1095_
timestamp 1607721120
transform 1 0 40664 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1068_
timestamp 1607721120
transform 1 0 39008 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_5_451
timestamp 1607721120
transform 1 0 42596 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_439
timestamp 1607721120
transform 1 0 41492 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0891_
timestamp 1607721120
transform 1 0 42228 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_469
timestamp 1607721120
transform 1 0 44252 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_459
timestamp 1607721120
transform 1 0 43332 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1075_
timestamp 1607721120
transform 1 0 43424 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_487
timestamp 1607721120
transform 1 0 45908 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_481
timestamp 1607721120
transform 1 0 45356 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1607721120
transform 1 0 46000 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1288_
timestamp 1607721120
transform 1 0 46092 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_5_520
timestamp 1607721120
transform 1 0 48944 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_508
timestamp 1607721120
transform 1 0 47840 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _1080_
timestamp 1607721120
transform 1 0 49220 0 1 4896
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_5_548
timestamp 1607721120
transform 1 0 51520 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_536
timestamp 1607721120
transform 1 0 50416 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_568
timestamp 1607721120
transform 1 0 53360 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_558
timestamp 1607721120
transform 1 0 52440 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_550
timestamp 1607721120
transform 1 0 51704 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1607721120
transform 1 0 51612 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1049_
timestamp 1607721120
transform 1 0 52532 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_591
timestamp 1607721120
transform 1 0 55476 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_580
timestamp 1607721120
transform 1 0 54464 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1082_
timestamp 1607721120
transform 1 0 54648 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_616
timestamp 1607721120
transform 1 0 57776 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_611
timestamp 1607721120
transform 1 0 57316 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_609
timestamp 1607721120
transform 1 0 57132 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_603
timestamp 1607721120
transform 1 0 56580 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1607721120
transform 1 0 57224 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0659_
timestamp 1607721120
transform 1 0 57408 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1289_
timestamp 1607721120
transform 1 0 58512 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_5_655
timestamp 1607721120
transform 1 0 61364 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_643
timestamp 1607721120
transform 1 0 60260 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1607721120
transform -1 0 62192 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_20
timestamp 1607721120
transform 1 0 2944 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1607721120
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1607721120
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_15
timestamp 1607721120
transform 1 0 2484 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1607721120
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1607721120
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1607721120
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1186_
timestamp 1607721120
transform 1 0 2668 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1173_
timestamp 1607721120
transform 1 0 2576 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_7_40
timestamp 1607721120
transform 1 0 4784 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_45
timestamp 1607721120
transform 1 0 5244 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_32
timestamp 1607721120
transform 1 0 4048 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1607721120
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1607721120
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1178_
timestamp 1607721120
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _1176_
timestamp 1607721120
transform 1 0 3680 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1607721120
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_52
timestamp 1607721120
transform 1 0 5888 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_66
timestamp 1607721120
transform 1 0 7176 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1607721120
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0932_
timestamp 1607721120
transform 1 0 6808 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _0928_
timestamp 1607721120
transform 1 0 5980 0 -1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1607721120
transform 1 0 8464 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_69
timestamp 1607721120
transform 1 0 7452 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1607721120
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_83
timestamp 1607721120
transform 1 0 8740 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0930_
timestamp 1607721120
transform 1 0 7912 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1607721120
transform 1 0 8188 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_106
timestamp 1607721120
transform 1 0 10856 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_105
timestamp 1607721120
transform 1 0 10764 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1607721120
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1607721120
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1308_
timestamp 1607721120
transform 1 0 11040 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__a211o_4  _0989_
timestamp 1607721120
transform 1 0 9568 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_7_132
timestamp 1607721120
transform 1 0 13248 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1607721120
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_127
timestamp 1607721120
transform 1 0 12788 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1607721120
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0890_
timestamp 1607721120
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0814_
timestamp 1607721120
transform 1 0 13524 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_158
timestamp 1607721120
transform 1 0 15640 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_150
timestamp 1607721120
transform 1 0 14904 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_144
timestamp 1607721120
transform 1 0 14352 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1607721120
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1607721120
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_139
timestamp 1607721120
transform 1 0 13892 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1607721120
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0974_
timestamp 1607721120
transform 1 0 14996 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0909_
timestamp 1607721120
transform 1 0 15456 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_7_175
timestamp 1607721120
transform 1 0 17204 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_163
timestamp 1607721120
transform 1 0 16100 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1312_
timestamp 1607721120
transform 1 0 16836 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__or3_4  _0978_
timestamp 1607721120
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_196
timestamp 1607721120
transform 1 0 19136 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_188
timestamp 1607721120
transform 1 0 18400 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_205
timestamp 1607721120
transform 1 0 19964 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_190
timestamp 1607721120
transform 1 0 18584 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1607721120
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_4  _0963_
timestamp 1607721120
transform 1 0 19320 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_4  _0907_
timestamp 1607721120
transform 1 0 19320 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0902_
timestamp 1607721120
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_228
timestamp 1607721120
transform 1 0 22080 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_211
timestamp 1607721120
transform 1 0 20516 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1607721120
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1607721120
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1607721120
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1607721120
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1185_
timestamp 1607721120
transform 1 0 21252 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_7_251
timestamp 1607721120
transform 1 0 24196 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_245
timestamp 1607721120
transform 1 0 23644 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_240
timestamp 1607721120
transform 1 0 23184 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_248
timestamp 1607721120
transform 1 0 23920 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1607721120
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0945_
timestamp 1607721120
transform 1 0 23092 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0898_
timestamp 1607721120
transform 1 0 23828 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_273
timestamp 1607721120
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp 1607721120
transform 1 0 25484 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1249_
timestamp 1607721120
transform 1 0 24932 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _0944_
timestamp 1607721120
transform 1 0 24656 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_7_296
timestamp 1607721120
transform 1 0 28336 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_290
timestamp 1607721120
transform 1 0 27784 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_278
timestamp 1607721120
transform 1 0 26680 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_293
timestamp 1607721120
transform 1 0 28060 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1607721120
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__a41o_4  _0957_
timestamp 1607721120
transform 1 0 26496 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _0824_
timestamp 1607721120
transform 1 0 27968 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_310
timestamp 1607721120
transform 1 0 29624 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_304
timestamp 1607721120
transform 1 0 29072 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_308
timestamp 1607721120
transform 1 0 29440 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1607721120
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1107_
timestamp 1607721120
transform 1 0 30176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0833_
timestamp 1607721120
transform 1 0 29256 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _0817_
timestamp 1607721120
transform 1 0 28796 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_7_334
timestamp 1607721120
transform 1 0 31832 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_328
timestamp 1607721120
transform 1 0 31280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1607721120
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1104_
timestamp 1607721120
transform 1 0 30728 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0841_
timestamp 1607721120
transform 1 0 32108 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_7_358
timestamp 1607721120
transform 1 0 34040 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_350
timestamp 1607721120
transform 1 0 33304 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_346
timestamp 1607721120
transform 1 0 32936 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_360
timestamp 1607721120
transform 1 0 34224 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_356
timestamp 1607721120
transform 1 0 33856 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_344
timestamp 1607721120
transform 1 0 32752 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0999_
timestamp 1607721120
transform 1 0 33396 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0834_
timestamp 1607721120
transform 1 0 34316 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_7_371
timestamp 1607721120
transform 1 0 35236 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_388
timestamp 1607721120
transform 1 0 36800 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_380
timestamp 1607721120
transform 1 0 36064 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_368
timestamp 1607721120
transform 1 0 34960 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1607721120
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1055_
timestamp 1607721120
transform 1 0 35972 0 1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _0853_
timestamp 1607721120
transform 1 0 34868 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0650_
timestamp 1607721120
transform 1 0 36432 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_409
timestamp 1607721120
transform 1 0 38732 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_401
timestamp 1607721120
transform 1 0 37996 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_406
timestamp 1607721120
transform 1 0 38456 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_398
timestamp 1607721120
transform 1 0 37720 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_396
timestamp 1607721120
transform 1 0 37536 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1607721120
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0854_
timestamp 1607721120
transform 1 0 38088 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_419
timestamp 1607721120
transform 1 0 39652 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_421
timestamp 1607721120
transform 1 0 39836 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1607721120
transform 1 0 40388 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1161_
timestamp 1607721120
transform 1 0 39008 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _1096_
timestamp 1607721120
transform 1 0 40572 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _1094_
timestamp 1607721120
transform 1 0 39192 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1024_
timestamp 1607721120
transform 1 0 40480 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_7_456
timestamp 1607721120
transform 1 0 43056 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_435
timestamp 1607721120
transform 1 0 41124 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_450
timestamp 1607721120
transform 1 0 42504 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_438
timestamp 1607721120
transform 1 0 41400 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1054_
timestamp 1607721120
transform 1 0 41860 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _0835_
timestamp 1607721120
transform 1 0 42136 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_472
timestamp 1607721120
transform 1 0 44528 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_468
timestamp 1607721120
transform 1 0 44160 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_473
timestamp 1607721120
transform 1 0 44620 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_463
timestamp 1607721120
transform 1 0 43700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_459
timestamp 1607721120
transform 1 0 43332 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1607721120
transform 1 0 43240 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1151_
timestamp 1607721120
transform 1 0 44620 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1073_
timestamp 1607721120
transform 1 0 43792 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_7_499
timestamp 1607721120
transform 1 0 47012 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_489
timestamp 1607721120
transform 1 0 46092 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_480
timestamp 1607721120
transform 1 0 45264 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_498
timestamp 1607721120
transform 1 0 46920 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_490
timestamp 1607721120
transform 1 0 46184 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1607721120
transform 1 0 46000 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1078_
timestamp 1607721120
transform 1 0 45356 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _1077_
timestamp 1607721120
transform 1 0 47012 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1062_
timestamp 1607721120
transform 1 0 46368 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_7_520
timestamp 1607721120
transform 1 0 48944 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_520
timestamp 1607721120
transform 1 0 48944 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_511
timestamp 1607721120
transform 1 0 48116 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1607721120
transform 1 0 48852 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_4  _1063_
timestamp 1607721120
transform 1 0 47748 0 1 5984
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_4  _1053_
timestamp 1607721120
transform 1 0 49220 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_7_541
timestamp 1607721120
transform 1 0 50876 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_532
timestamp 1607721120
transform 1 0 50048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_544
timestamp 1607721120
transform 1 0 51152 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_532
timestamp 1607721120
transform 1 0 50048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _1076_
timestamp 1607721120
transform 1 0 50232 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1064_
timestamp 1607721120
transform 1 0 51520 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_7_556
timestamp 1607721120
transform 1 0 52256 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_550
timestamp 1607721120
transform 1 0 51704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_555
timestamp 1607721120
transform 1 0 52164 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1607721120
transform 1 0 51612 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1058_
timestamp 1607721120
transform 1 0 51888 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _1052_
timestamp 1607721120
transform 1 0 52900 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _1050_
timestamp 1607721120
transform 1 0 52992 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_7_593
timestamp 1607721120
transform 1 0 55660 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_573
timestamp 1607721120
transform 1 0 53820 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_581
timestamp 1607721120
transform 1 0 54556 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_572
timestamp 1607721120
transform 1 0 53728 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1607721120
transform 1 0 54464 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1066_
timestamp 1607721120
transform 1 0 54556 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _1065_
timestamp 1607721120
transform 1 0 55292 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_611
timestamp 1607721120
transform 1 0 57316 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_609
timestamp 1607721120
transform 1 0 57132 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_605
timestamp 1607721120
transform 1 0 56764 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_601
timestamp 1607721120
transform 1 0 56396 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1607721120
transform 1 0 57224 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1069_
timestamp 1607721120
transform 1 0 57132 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_7_633
timestamp 1607721120
transform 1 0 59340 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_637
timestamp 1607721120
transform 1 0 59708 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_625
timestamp 1607721120
transform 1 0 58604 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _1072_
timestamp 1607721120
transform 1 0 58052 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_7_653
timestamp 1607721120
transform 1 0 61180 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_649
timestamp 1607721120
transform 1 0 60812 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1607721120
transform 1 0 60076 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1607721120
transform -1 0 62192 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1607721120
transform -1 0 62192 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1071_
timestamp 1607721120
transform 1 0 60168 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _1056_
timestamp 1607721120
transform 1 0 60076 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_19
timestamp 1607721120
transform 1 0 2852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1607721120
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1607721120
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1607721120
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1184_
timestamp 1607721120
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_23
timestamp 1607721120
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1607721120
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1250_
timestamp 1607721120
transform 1 0 4048 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_8_66
timestamp 1607721120
transform 1 0 7176 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_51
timestamp 1607721120
transform 1 0 5796 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1177_
timestamp 1607721120
transform 1 0 6532 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_8_84
timestamp 1607721120
transform 1 0 8832 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_74
timestamp 1607721120
transform 1 0 7912 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _0987_
timestamp 1607721120
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_108
timestamp 1607721120
transform 1 0 11040 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1607721120
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a21boi_4  _0988_
timestamp 1607721120
transform 1 0 9660 0 -1 7072
box -38 -48 1418 592
use sky130_fd_sc_hd__fill_1  FILLER_8_137
timestamp 1607721120
transform 1 0 13708 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_129
timestamp 1607721120
transform 1 0 12972 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_4  _0986_
timestamp 1607721120
transform 1 0 11776 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_8_154
timestamp 1607721120
transform 1 0 15272 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_145
timestamp 1607721120
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1607721120
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0995_
timestamp 1607721120
transform 1 0 13800 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_8_181
timestamp 1607721120
transform 1 0 17756 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1304_
timestamp 1607721120
transform 1 0 16008 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_8_205
timestamp 1607721120
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_189
timestamp 1607721120
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0967_
timestamp 1607721120
transform 1 0 18676 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_8_224
timestamp 1607721120
transform 1 0 21712 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1607721120
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1607721120
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _0973_
timestamp 1607721120
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_243
timestamp 1607721120
transform 1 0 23460 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0847_
timestamp 1607721120
transform 1 0 22816 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_8_267
timestamp 1607721120
transform 1 0 25668 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _1180_
timestamp 1607721120
transform 1 0 24564 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_276
timestamp 1607721120
transform 1 0 26496 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1607721120
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _0955_
timestamp 1607721120
transform 1 0 26772 0 -1 7072
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_8  FILLER_8_316
timestamp 1607721120
transform 1 0 30176 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_309
timestamp 1607721120
transform 1 0 29532 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_301
timestamp 1607721120
transform 1 0 28796 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0882_
timestamp 1607721120
transform 1 0 29808 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_337
timestamp 1607721120
transform 1 0 32108 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_328
timestamp 1607721120
transform 1 0 31280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1607721120
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0820_
timestamp 1607721120
transform 1 0 30912 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_364
timestamp 1607721120
transform 1 0 34592 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_347
timestamp 1607721120
transform 1 0 33028 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _1183_
timestamp 1607721120
transform 1 0 33764 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0837_
timestamp 1607721120
transform 1 0 32660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_4  _1007_
timestamp 1607721120
transform 1 0 35328 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_8_401
timestamp 1607721120
transform 1 0 37996 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_389
timestamp 1607721120
transform 1 0 36892 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1607721120
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1045_
timestamp 1607721120
transform 1 0 38732 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1607721120
transform 1 0 37720 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_433
timestamp 1607721120
transform 1 0 40940 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_416
timestamp 1607721120
transform 1 0 39376 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1047_
timestamp 1607721120
transform 1 0 40112 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_450
timestamp 1607721120
transform 1 0 42504 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1025_
timestamp 1607721120
transform 1 0 41676 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_471
timestamp 1607721120
transform 1 0 44436 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1607721120
transform 1 0 43240 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1028_
timestamp 1607721120
transform 1 0 45172 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _1016_
timestamp 1607721120
transform 1 0 43332 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_488
timestamp 1607721120
transform 1 0 46000 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _1181_
timestamp 1607721120
transform 1 0 46736 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_517
timestamp 1607721120
transform 1 0 48668 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_505
timestamp 1607721120
transform 1 0 47564 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1607721120
transform 1 0 48852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1149_
timestamp 1607721120
transform 1 0 48944 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_8_539
timestamp 1607721120
transform 1 0 50692 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_527
timestamp 1607721120
transform 1 0 49588 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _1155_
timestamp 1607721120
transform 1 0 51060 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_8_550
timestamp 1607721120
transform 1 0 51704 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1067_
timestamp 1607721120
transform 1 0 52440 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_8_590
timestamp 1607721120
transform 1 0 55384 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_581
timestamp 1607721120
transform 1 0 54556 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_572
timestamp 1607721120
transform 1 0 53728 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1607721120
transform 1 0 54464 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1051_
timestamp 1607721120
transform 1 0 54740 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_8_611
timestamp 1607721120
transform 1 0 57316 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1059_
timestamp 1607721120
transform 1 0 56120 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_8_633
timestamp 1607721120
transform 1 0 59340 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1061_
timestamp 1607721120
transform 1 0 58052 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_8_649
timestamp 1607721120
transform 1 0 60812 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1607721120
transform 1 0 60076 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1607721120
transform -1 0 62192 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1157_
timestamp 1607721120
transform 1 0 60168 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1607721120
transform 1 0 2484 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1607721120
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1607721120
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1251_
timestamp 1607721120
transform 1 0 2852 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_9_38
timestamp 1607721120
transform 1 0 4600 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1607721120
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_53
timestamp 1607721120
transform 1 0 5980 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1607721120
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1175_
timestamp 1607721120
transform 1 0 5336 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_74
timestamp 1607721120
transform 1 0 7912 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1302_
timestamp 1607721120
transform 1 0 8280 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_9_114
timestamp 1607721120
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_97
timestamp 1607721120
transform 1 0 10028 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0982_
timestamp 1607721120
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_137
timestamp 1607721120
transform 1 0 13708 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1607721120
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0983_
timestamp 1607721120
transform 1 0 12420 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_9_152
timestamp 1607721120
transform 1 0 15088 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1121_
timestamp 1607721120
transform 1 0 14444 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_9_175
timestamp 1607721120
transform 1 0 17204 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_165
timestamp 1607721120
transform 1 0 16284 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_160
timestamp 1607721120
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 16008 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _0975_
timestamp 1607721120
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_188
timestamp 1607721120
transform 1 0 18400 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1607721120
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1607721120
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1306_
timestamp 1607721120
transform 1 0 18492 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_9_228
timestamp 1607721120
transform 1 0 22080 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_208
timestamp 1607721120
transform 1 0 20240 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _0965_
timestamp 1607721120
transform 1 0 20976 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_245
timestamp 1607721120
transform 1 0 23644 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_240
timestamp 1607721120
transform 1 0 23184 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1607721120
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1179_
timestamp 1607721120
transform 1 0 24196 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_9_270
timestamp 1607721120
transform 1 0 25944 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_258
timestamp 1607721120
transform 1 0 24840 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0958_
timestamp 1607721120
transform 1 0 25576 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_292
timestamp 1607721120
transform 1 0 27968 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1607721120
transform 1 0 26680 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0956_
timestamp 1607721120
transform 1 0 26864 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_313
timestamp 1607721120
transform 1 0 29900 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_304
timestamp 1607721120
transform 1 0 29072 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1607721120
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0950_
timestamp 1607721120
transform 1 0 29256 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1607721120
transform 1 0 32108 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_325
timestamp 1607721120
transform 1 0 31004 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0839_
timestamp 1607721120
transform 1 0 31740 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0838_
timestamp 1607721120
transform 1 0 30636 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_358
timestamp 1607721120
transform 1 0 34040 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1145_
timestamp 1607721120
transform 1 0 33212 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_371
timestamp 1607721120
transform 1 0 35236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_367
timestamp 1607721120
transform 1 0 34868 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1607721120
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a41oi_4  _1005_
timestamp 1607721120
transform 1 0 35328 0 1 7072
box -38 -48 2062 592
use sky130_fd_sc_hd__decap_6  FILLER_9_406
timestamp 1607721120
transform 1 0 38456 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_394
timestamp 1607721120
transform 1 0 37352 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_428
timestamp 1607721120
transform 1 0 40480 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_419
timestamp 1607721120
transform 1 0 39652 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1607721120
transform 1 0 40388 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1012_
timestamp 1607721120
transform 1 0 39008 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_9_448
timestamp 1607721120
transform 1 0 42320 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_434
timestamp 1607721120
transform 1 0 41032 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_4  _1013_
timestamp 1607721120
transform 1 0 41124 0 1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _0906_
timestamp 1607721120
transform 1 0 43056 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_460
timestamp 1607721120
transform 1 0 43424 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1015_
timestamp 1607721120
transform 1 0 44160 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_501
timestamp 1607721120
transform 1 0 47196 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_480
timestamp 1607721120
transform 1 0 45264 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1607721120
transform 1 0 46000 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1027_
timestamp 1607721120
transform 1 0 46092 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_521
timestamp 1607721120
transform 1 0 49036 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_513
timestamp 1607721120
transform 1 0 48300 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0868_
timestamp 1607721120
transform 1 0 48668 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_541
timestamp 1607721120
transform 1 0 50876 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_533
timestamp 1607721120
transform 1 0 50140 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1039_
timestamp 1607721120
transform 1 0 50508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_550
timestamp 1607721120
transform 1 0 51704 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1607721120
transform 1 0 51612 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1290_
timestamp 1607721120
transform 1 0 52256 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_9_587
timestamp 1607721120
transform 1 0 55108 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_575
timestamp 1607721120
transform 1 0 54004 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_4  _1037_
timestamp 1607721120
transform 1 0 55660 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_615
timestamp 1607721120
transform 1 0 57684 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_602
timestamp 1607721120
transform 1 0 56488 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1607721120
transform 1 0 57224 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0864_
timestamp 1607721120
transform 1 0 57316 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_623
timestamp 1607721120
transform 1 0 58420 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1291_
timestamp 1607721120
transform 1 0 58512 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_9_655
timestamp 1607721120
transform 1 0 61364 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_643
timestamp 1607721120
transform 1 0 60260 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1607721120
transform -1 0 62192 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1607721120
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1607721120
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _1174_
timestamp 1607721120
transform 1 0 2116 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1607721120
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_23
timestamp 1607721120
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1607721120
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1170_
timestamp 1607721120
transform 1 0 4232 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_58
timestamp 1607721120
transform 1 0 6440 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_46
timestamp 1607721120
transform 1 0 5336 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1607721120
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_76
timestamp 1607721120
transform 1 0 8096 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_70
timestamp 1607721120
transform 1 0 7544 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0981_
timestamp 1607721120
transform 1 0 8188 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_10_107
timestamp 1607721120
transform 1 0 10948 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1607721120
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0991_
timestamp 1607721120
transform 1 0 9660 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_10_131
timestamp 1607721120
transform 1 0 13156 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_115
timestamp 1607721120
transform 1 0 11684 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_wb_clk_i
timestamp 1607721120
transform 1 0 11776 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _0985_
timestamp 1607721120
transform 1 0 12052 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_145
timestamp 1607721120
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_139
timestamp 1607721120
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1607721120
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1123_
timestamp 1607721120
transform 1 0 15272 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0970_
timestamp 1607721120
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_182
timestamp 1607721120
transform 1 0 17848 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_169
timestamp 1607721120
transform 1 0 16652 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_161
timestamp 1607721120
transform 1 0 15916 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _0977_
timestamp 1607721120
transform 1 0 16744 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _0966_
timestamp 1607721120
transform 1 0 18952 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_222
timestamp 1607721120
transform 1 0 21528 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_206
timestamp 1607721120
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1607721120
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0962_
timestamp 1607721120
transform 1 0 20884 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_10_243
timestamp 1607721120
transform 1 0 23460 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_4  _0954_
timestamp 1607721120
transform 1 0 22264 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_10_267
timestamp 1607721120
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_255
timestamp 1607721120
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_293
timestamp 1607721120
transform 1 0 28060 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_276
timestamp 1607721120
transform 1 0 26496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1607721120
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0961_
timestamp 1607721120
transform 1 0 26772 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_10_310
timestamp 1607721120
transform 1 0 29624 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1109_
timestamp 1607721120
transform 1 0 30360 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _0960_
timestamp 1607721120
transform 1 0 28796 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_337
timestamp 1607721120
transform 1 0 32108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_335
timestamp 1607721120
transform 1 0 31924 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_327
timestamp 1607721120
transform 1 0 31188 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1607721120
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0844_
timestamp 1607721120
transform 1 0 32476 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_10_348
timestamp 1607721120
transform 1 0 33120 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1011_
timestamp 1607721120
transform 1 0 33856 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_10_387
timestamp 1607721120
transform 1 0 36708 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_370
timestamp 1607721120
transform 1 0 35144 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1010_
timestamp 1607721120
transform 1 0 35880 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_410
timestamp 1607721120
transform 1 0 38824 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_402
timestamp 1607721120
transform 1 0 38088 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_395
timestamp 1607721120
transform 1 0 37444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1607721120
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0888_
timestamp 1607721120
transform 1 0 37720 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_419
timestamp 1607721120
transform 1 0 39652 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1135_
timestamp 1607721120
transform 1 0 39008 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_4  _1046_
timestamp 1607721120
transform 1 0 40388 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_456
timestamp 1607721120
transform 1 0 43056 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_448
timestamp 1607721120
transform 1 0 42320 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_436
timestamp 1607721120
transform 1 0 41216 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1008_
timestamp 1607721120
transform 1 0 41952 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_476
timestamp 1607721120
transform 1 0 44896 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_468
timestamp 1607721120
transform 1 0 44160 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1607721120
transform 1 0 43240 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1296_
timestamp 1607721120
transform 1 0 45080 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1023_
timestamp 1607721120
transform 1 0 43332 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_497
timestamp 1607721120
transform 1 0 46828 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_520
timestamp 1607721120
transform 1 0 48944 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_517
timestamp 1607721120
transform 1 0 48668 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_509
timestamp 1607721120
transform 1 0 47932 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1607721120
transform 1 0 48852 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1020_
timestamp 1607721120
transform 1 0 47564 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_532
timestamp 1607721120
transform 1 0 50048 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1030_
timestamp 1607721120
transform 1 0 50600 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_10_563
timestamp 1607721120
transform 1 0 52900 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_551
timestamp 1607721120
transform 1 0 51796 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _1147_
timestamp 1607721120
transform 1 0 53084 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_10_592
timestamp 1607721120
transform 1 0 55568 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_581
timestamp 1607721120
transform 1 0 54556 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_572
timestamp 1607721120
transform 1 0 53728 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1607721120
transform 1 0 54464 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1032_
timestamp 1607721120
transform 1 0 54740 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_614
timestamp 1607721120
transform 1 0 57592 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _1042_
timestamp 1607721120
transform 1 0 56304 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_10_639
timestamp 1607721120
transform 1 0 59892 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_631
timestamp 1607721120
transform 1 0 59156 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1060_
timestamp 1607721120
transform 1 0 58328 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_649
timestamp 1607721120
transform 1 0 60812 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1607721120
transform 1 0 60076 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1607721120
transform -1 0 62192 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1159_
timestamp 1607721120
transform 1 0 60168 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_11_11
timestamp 1607721120
transform 1 0 2116 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1607721120
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1607721120
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1607721120
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1252_
timestamp 1607721120
transform 1 0 2852 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1182_
timestamp 1607721120
transform 1 0 1840 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_38
timestamp 1607721120
transform 1 0 4600 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1607721120
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_58
timestamp 1607721120
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_50
timestamp 1607721120
transform 1 0 5704 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1607721120
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1164_
timestamp 1607721120
transform 1 0 5336 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_74
timestamp 1607721120
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1301_
timestamp 1607721120
transform 1 0 8096 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_11_112
timestamp 1607721120
transform 1 0 11408 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_95
timestamp 1607721120
transform 1 0 9844 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _0996_
timestamp 1607721120
transform 1 0 10580 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_123
timestamp 1607721120
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1607721120
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1607721120
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _0980_
timestamp 1607721120
transform 1 0 12696 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_11_158
timestamp 1607721120
transform 1 0 15640 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_150
timestamp 1607721120
transform 1 0 14904 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_139
timestamp 1607721120
transform 1 0 13892 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1607721120
transform 1 0 14628 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_180
timestamp 1607721120
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_168
timestamp 1607721120
transform 1 0 16560 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0976_
timestamp 1607721120
transform 1 0 15916 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_11_196
timestamp 1607721120
transform 1 0 19136 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_188
timestamp 1607721120
transform 1 0 18400 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_184
timestamp 1607721120
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1607721120
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0969_
timestamp 1607721120
transform 1 0 19872 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_4  _0964_
timestamp 1607721120
transform 1 0 18492 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_11_220
timestamp 1607721120
transform 1 0 21344 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0968_
timestamp 1607721120
transform 1 0 22080 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_11_249
timestamp 1607721120
transform 1 0 24012 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_243
timestamp 1607721120
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_235
timestamp 1607721120
transform 1 0 22724 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1607721120
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0848_
timestamp 1607721120
transform 1 0 23644 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_268
timestamp 1607721120
transform 1 0 25760 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_257
timestamp 1607721120
transform 1 0 24748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0865_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 24932 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_289
timestamp 1607721120
transform 1 0 27692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _0959_
timestamp 1607721120
transform 1 0 26496 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1607721120
transform 1 0 30268 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_306
timestamp 1607721120
transform 1 0 29256 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_301
timestamp 1607721120
transform 1 0 28796 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1607721120
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1111_
timestamp 1607721120
transform 1 0 29624 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_11_341
timestamp 1607721120
transform 1 0 32476 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_333
timestamp 1607721120
transform 1 0 31740 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_329
timestamp 1607721120
transform 1 0 31372 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1139_
timestamp 1607721120
transform 1 0 31832 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_11_358
timestamp 1607721120
transform 1 0 34040 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1127_
timestamp 1607721120
transform 1 0 33212 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_380
timestamp 1607721120
transform 1 0 36064 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1607721120
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1143_
timestamp 1607721120
transform 1 0 36800 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1009_
timestamp 1607721120
transform 1 0 34868 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_11_407
timestamp 1607721120
transform 1 0 38548 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_395
timestamp 1607721120
transform 1 0 37444 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0845_
timestamp 1607721120
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_432
timestamp 1607721120
transform 1 0 40848 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_419
timestamp 1607721120
transform 1 0 39652 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1607721120
transform 1 0 40388 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0920_
timestamp 1607721120
transform 1 0 39284 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0904_
timestamp 1607721120
transform 1 0 40480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_454
timestamp 1607721120
transform 1 0 42872 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1017_
timestamp 1607721120
transform 1 0 41584 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_11_476
timestamp 1607721120
transform 1 0 44896 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1022_
timestamp 1607721120
transform 1 0 43608 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_11_502
timestamp 1607721120
transform 1 0 47288 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_487
timestamp 1607721120
transform 1 0 45908 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_wb_clk_i
timestamp 1607721120
transform 1 0 45632 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1607721120
transform 1 0 46000 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1004_
timestamp 1607721120
transform 1 0 46092 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_11_517
timestamp 1607721120
transform 1 0 48668 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1014_
timestamp 1607721120
transform 1 0 48024 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_11_541
timestamp 1607721120
transform 1 0 50876 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_533
timestamp 1607721120
transform 1 0 50140 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_529
timestamp 1607721120
transform 1 0 49772 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1026_
timestamp 1607721120
transform 1 0 50232 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_11_558
timestamp 1607721120
transform 1 0 52440 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_550
timestamp 1607721120
transform 1 0 51704 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1607721120
transform 1 0 51612 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1048_
timestamp 1607721120
transform 1 0 52624 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  FILLER_11_582
timestamp 1607721120
transform 1 0 54648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_574
timestamp 1607721120
transform 1 0 53912 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_4  _1036_
timestamp 1607721120
transform 1 0 54924 0 1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_11_611
timestamp 1607721120
transform 1 0 57316 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_598
timestamp 1607721120
transform 1 0 56120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1607721120
transform 1 0 57224 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_639
timestamp 1607721120
transform 1 0 59892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_623
timestamp 1607721120
transform 1 0 58420 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a21boi_4  _1038_
timestamp 1607721120
transform 1 0 58512 0 1 8160
box -38 -48 1418 592
use sky130_fd_sc_hd__fill_2  FILLER_11_659
timestamp 1607721120
transform 1 0 61732 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_651
timestamp 1607721120
transform 1 0 60996 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1607721120
transform -1 0 62192 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1607721120
transform 1 0 1380 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1607721120
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _1172_
timestamp 1607721120
transform 1 0 2116 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_38
timestamp 1607721120
transform 1 0 4600 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_32
timestamp 1607721120
transform 1 0 4048 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1607721120
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1607721120
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1166_
timestamp 1607721120
transform 1 0 4692 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_63
timestamp 1607721120
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_51
timestamp 1607721120
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_84
timestamp 1607721120
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_75
timestamp 1607721120
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0992_
timestamp 1607721120
transform 1 0 8188 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_107
timestamp 1607721120
transform 1 0 10948 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1607721120
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0994_
timestamp 1607721120
transform 1 0 9660 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_12_129
timestamp 1607721120
transform 1 0 12972 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0998_
timestamp 1607721120
transform 1 0 11684 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_4  _0984_
timestamp 1607721120
transform 1 0 13708 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_154
timestamp 1607721120
transform 1 0 15272 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1607721120
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_144
timestamp 1607721120
transform 1 0 14352 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1607721120
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_174
timestamp 1607721120
transform 1 0 17112 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_165
timestamp 1607721120
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_wb_clk_i
timestamp 1607721120
transform 1 0 16008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1119_
timestamp 1607721120
transform 1 0 16468 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0971_
timestamp 1607721120
transform 1 0 17848 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_189
timestamp 1607721120
transform 1 0 18492 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0949_
timestamp 1607721120
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_206
timestamp 1607721120
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1607721120
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0972_
timestamp 1607721120
transform 1 0 20884 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_12_246
timestamp 1607721120
transform 1 0 23736 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_229
timestamp 1607721120
transform 1 0 22172 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _0952_
timestamp 1607721120
transform 1 0 22908 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_272
timestamp 1607721120
transform 1 0 26128 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_260
timestamp 1607721120
transform 1 0 25024 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_254
timestamp 1607721120
transform 1 0 24472 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1607721120
transform 1 0 24748 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_276
timestamp 1607721120
transform 1 0 26496 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1607721120
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1307_
timestamp 1607721120
transform 1 0 27048 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_12_318
timestamp 1607721120
transform 1 0 30360 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_313
timestamp 1607721120
transform 1 0 29900 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_301
timestamp 1607721120
transform 1 0 28796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0886_
timestamp 1607721120
transform 1 0 29992 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_340
timestamp 1607721120
transform 1 0 32384 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_333
timestamp 1607721120
transform 1 0 31740 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_325
timestamp 1607721120
transform 1 0 31004 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1607721120
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0901_
timestamp 1607721120
transform 1 0 30636 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1607721120
transform 1 0 32108 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1299_
timestamp 1607721120
transform 1 0 33120 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_12_387
timestamp 1607721120
transform 1 0 36708 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_367
timestamp 1607721120
transform 1 0 34868 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _1144_
timestamp 1607721120
transform 1 0 35604 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_405
timestamp 1607721120
transform 1 0 38364 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_395
timestamp 1607721120
transform 1 0 37444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1607721120
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1129_
timestamp 1607721120
transform 1 0 37720 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_428
timestamp 1607721120
transform 1 0 40480 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_417
timestamp 1607721120
transform 1 0 39468 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _1018_
timestamp 1607721120
transform 1 0 39836 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_12_455
timestamp 1607721120
transform 1 0 42964 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_443
timestamp 1607721120
transform 1 0 41860 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _1131_
timestamp 1607721120
transform 1 0 41216 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_12_465
timestamp 1607721120
transform 1 0 43884 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_459
timestamp 1607721120
transform 1 0 43332 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1607721120
transform 1 0 43240 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1019_
timestamp 1607721120
transform 1 0 43976 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_499
timestamp 1607721120
transform 1 0 47012 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_482
timestamp 1607721120
transform 1 0 45448 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _1003_
timestamp 1607721120
transform 1 0 46184 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_524
timestamp 1607721120
transform 1 0 49312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_520
timestamp 1607721120
transform 1 0 48944 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_518
timestamp 1607721120
transform 1 0 48760 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_510
timestamp 1607721120
transform 1 0 48024 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_wb_clk_i
timestamp 1607721120
transform 1 0 47748 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1607721120
transform 1 0 48852 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1034_
timestamp 1607721120
transform 1 0 49404 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_532
timestamp 1607721120
transform 1 0 50048 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _1033_
timestamp 1607721120
transform 1 0 50784 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_12_554
timestamp 1607721120
transform 1 0 52072 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1000_
timestamp 1607721120
transform 1 0 52808 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_589
timestamp 1607721120
transform 1 0 55292 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_581
timestamp 1607721120
transform 1 0 54556 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_579
timestamp 1607721120
transform 1 0 54372 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_571
timestamp 1607721120
transform 1 0 53636 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1607721120
transform 1 0 54464 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1041_
timestamp 1607721120
transform 1 0 54648 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_611
timestamp 1607721120
transform 1 0 57316 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1044_
timestamp 1607721120
transform 1 0 56028 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_12_633
timestamp 1607721120
transform 1 0 59340 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1040_
timestamp 1607721120
transform 1 0 58052 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_12_649
timestamp 1607721120
transform 1 0 60812 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1607721120
transform 1 0 60076 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1607721120
transform -1 0 62192 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1043_
timestamp 1607721120
transform 1 0 60168 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1607721120
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1607721120
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_19
timestamp 1607721120
transform 1 0 2852 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 1607721120
transform 1 0 2484 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1607721120
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1607721120
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1607721120
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1253_
timestamp 1607721120
transform 1 0 2944 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1607721120
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1607721120
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1607721120
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1254_
timestamp 1607721120
transform 1 0 4048 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_14_66
timestamp 1607721120
transform 1 0 7176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_51
timestamp 1607721120
transform 1 0 5796 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1607721120
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1607721120
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1607721120
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1168_
timestamp 1607721120
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0810_
timestamp 1607721120
transform 1 0 6532 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1607721120
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_78
timestamp 1607721120
transform 1 0 8280 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_74
timestamp 1607721120
transform 1 0 7912 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1300_
timestamp 1607721120
transform 1 0 8648 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_14_111
timestamp 1607721120
transform 1 0 11316 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_103
timestamp 1607721120
transform 1 0 10580 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1607721120
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1607721120
transform 1 0 11500 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_101
timestamp 1607721120
transform 1 0 10396 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1607721120
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0990_
timestamp 1607721120
transform 1 0 9936 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0798_
timestamp 1607721120
transform 1 0 11408 0 -1 10336
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _0768_
timestamp 1607721120
transform 1 0 11132 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_126
timestamp 1607721120
transform 1 0 12696 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1607721120
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1607721120
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1303_
timestamp 1607721120
transform 1 0 12420 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__or4_4  _0948_
timestamp 1607721120
transform 1 0 13432 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1607721120
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_143
timestamp 1607721120
transform 1 0 14260 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_142
timestamp 1607721120
transform 1 0 14168 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1607721120
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1124_
timestamp 1607721120
transform 1 0 14904 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _1122_
timestamp 1607721120
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_178
timestamp 1607721120
transform 1 0 17480 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1607721120
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_175
timestamp 1607721120
transform 1 0 17204 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_170
timestamp 1607721120
transform 1 0 16744 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_162
timestamp 1607721120
transform 1 0 16008 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _1117_
timestamp 1607721120
transform 1 0 17848 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0860_
timestamp 1607721120
transform 1 0 16836 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_189
timestamp 1607721120
transform 1 0 18492 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_194
timestamp 1607721120
transform 1 0 18952 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_184
timestamp 1607721120
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1607721120
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1305_
timestamp 1607721120
transform 1 0 19688 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1113_
timestamp 1607721120
transform 1 0 18308 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _0953_
timestamp 1607721120
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_221
timestamp 1607721120
transform 1 0 21436 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_215
timestamp 1607721120
transform 1 0 20884 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_206
timestamp 1607721120
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_221
timestamp 1607721120
transform 1 0 21436 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1607721120
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0747_
timestamp 1607721120
transform 1 0 21068 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_248
timestamp 1607721120
transform 1 0 23920 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_248
timestamp 1607721120
transform 1 0 23920 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_236
timestamp 1607721120
transform 1 0 22816 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1607721120
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1317_
timestamp 1607721120
transform 1 0 22172 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1115_
timestamp 1607721120
transform 1 0 22172 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1607721120
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_267
timestamp 1607721120
transform 1 0 25668 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_270
timestamp 1607721120
transform 1 0 25944 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_260
timestamp 1607721120
transform 1 0 25024 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0867_
timestamp 1607721120
transform 1 0 25024 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0862_
timestamp 1607721120
transform 1 0 25300 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_14_293
timestamp 1607721120
transform 1 0 28060 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_295
timestamp 1607721120
transform 1 0 28244 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1607721120
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_4  _0871_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 26496 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__a32o_4  _0866_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 26680 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_14_308
timestamp 1607721120
transform 1 0 29440 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_313
timestamp 1607721120
transform 1 0 29900 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_303
timestamp 1607721120
transform 1 0 28980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1607721120
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1236_
timestamp 1607721120
transform 1 0 29256 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0946_
timestamp 1607721120
transform 1 0 30176 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _0858_
timestamp 1607721120
transform 1 0 28796 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_14_337
timestamp 1607721120
transform 1 0 32108 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_332
timestamp 1607721120
transform 1 0 31648 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_320
timestamp 1607721120
transform 1 0 30544 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_321
timestamp 1607721120
transform 1 0 30636 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607721120
transform 1 0 30728 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1607721120
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1141_
timestamp 1607721120
transform 1 0 32200 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0918_
timestamp 1607721120
transform 1 0 32568 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_345
timestamp 1607721120
transform 1 0 32844 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_358
timestamp 1607721120
transform 1 0 34040 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1265_
timestamp 1607721120
transform 1 0 33580 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _1142_
timestamp 1607721120
transform 1 0 32936 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_387
timestamp 1607721120
transform 1 0 36708 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_372
timestamp 1607721120
transform 1 0 35328 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_379
timestamp 1607721120
transform 1 0 35972 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1607721120
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1202_
timestamp 1607721120
transform 1 0 36064 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1137_
timestamp 1607721120
transform 1 0 36708 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _1006_
timestamp 1607721120
transform 1 0 34868 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_402
timestamp 1607721120
transform 1 0 38088 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_395
timestamp 1607721120
transform 1 0 37444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_406
timestamp 1607721120
transform 1 0 38456 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_394
timestamp 1607721120
transform 1 0 37352 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1607721120
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0951_
timestamp 1607721120
transform 1 0 37720 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_428
timestamp 1607721120
transform 1 0 40480 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_414
timestamp 1607721120
transform 1 0 39192 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_428
timestamp 1607721120
transform 1 0 40480 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_419
timestamp 1607721120
transform 1 0 39652 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1607721120
transform 1 0 40388 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1136_
timestamp 1607721120
transform 1 0 39376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _1133_
timestamp 1607721120
transform 1 0 39008 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_456
timestamp 1607721120
transform 1 0 43056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_448
timestamp 1607721120
transform 1 0 42320 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_439
timestamp 1607721120
transform 1 0 41492 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_wb_clk_i
timestamp 1607721120
transform 1 0 41216 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1298_
timestamp 1607721120
transform 1 0 41768 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _1132_
timestamp 1607721120
transform 1 0 41216 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_467
timestamp 1607721120
transform 1 0 44068 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_459
timestamp 1607721120
transform 1 0 43332 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_478
timestamp 1607721120
transform 1 0 45080 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_461
timestamp 1607721120
transform 1 0 43516 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1607721120
transform 1 0 43240 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1297_
timestamp 1607721120
transform 1 0 44344 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__or4_4  _1001_
timestamp 1607721120
transform 1 0 44252 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1607721120
transform 1 0 47196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_489
timestamp 1607721120
transform 1 0 46092 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_498
timestamp 1607721120
transform 1 0 46920 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_486
timestamp 1607721120
transform 1 0 45816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1607721120
transform 1 0 46000 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1002_
timestamp 1607721120
transform 1 0 46092 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0701_
timestamp 1607721120
transform 1 0 46828 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_513
timestamp 1607721120
transform 1 0 48300 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_524
timestamp 1607721120
transform 1 0 49312 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_513
timestamp 1607721120
transform 1 0 48300 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_wb_clk_i
timestamp 1607721120
transform 1 0 49036 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1607721120
transform 1 0 48852 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1150_
timestamp 1607721120
transform 1 0 48944 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _1021_
timestamp 1607721120
transform 1 0 47656 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_14_544
timestamp 1607721120
transform 1 0 51152 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_532
timestamp 1607721120
transform 1 0 50048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_541
timestamp 1607721120
transform 1 0 50876 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_528
timestamp 1607721120
transform 1 0 49680 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1295_
timestamp 1607721120
transform 1 0 51520 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _1035_
timestamp 1607721120
transform 1 0 49772 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_567
timestamp 1607721120
transform 1 0 53268 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_558
timestamp 1607721120
transform 1 0 52440 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_550
timestamp 1607721120
transform 1 0 51704 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1607721120
transform 1 0 51612 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1292_
timestamp 1607721120
transform 1 0 52624 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_14_586
timestamp 1607721120
transform 1 0 55016 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_581
timestamp 1607721120
transform 1 0 54556 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_579
timestamp 1607721120
transform 1 0 54372 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_587
timestamp 1607721120
transform 1 0 55108 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_579
timestamp 1607721120
transform 1 0 54372 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1607721120
transform 1 0 54464 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1031_
timestamp 1607721120
transform 1 0 55200 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0723_
timestamp 1607721120
transform 1 0 54648 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_606
timestamp 1607721120
transform 1 0 56856 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_611
timestamp 1607721120
transform 1 0 57316 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_607
timestamp 1607721120
transform 1 0 56948 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_595
timestamp 1607721120
transform 1 0 55844 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1607721120
transform 1 0 57224 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1294_
timestamp 1607721120
transform 1 0 57592 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _1158_
timestamp 1607721120
transform 1 0 55752 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_633
timestamp 1607721120
transform 1 0 59340 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_638
timestamp 1607721120
transform 1 0 59800 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1293_
timestamp 1607721120
transform 1 0 58052 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_14_660
timestamp 1607721120
transform 1 0 61824 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_654
timestamp 1607721120
transform 1 0 61272 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_642
timestamp 1607721120
transform 1 0 60168 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_658
timestamp 1607721120
transform 1 0 61640 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_650
timestamp 1607721120
transform 1 0 60904 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1607721120
transform 1 0 60076 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1607721120
transform -1 0 62192 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1607721120
transform -1 0 62192 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_15
timestamp 1607721120
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1607721120
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1607721120
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1233_
timestamp 1607721120
transform 1 0 2668 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_15_24
timestamp 1607721120
transform 1 0 3312 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1255_
timestamp 1607721120
transform 1 0 4048 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1607721120
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1607721120
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1607721120
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0801_
timestamp 1607721120
transform 1 0 6808 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_15_87
timestamp 1607721120
transform 1 0 9108 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_81
timestamp 1607721120
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1607721120
transform 1 0 7452 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0791_
timestamp 1607721120
transform 1 0 8740 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_114
timestamp 1607721120
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_99
timestamp 1607721120
transform 1 0 10212 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _0797_
timestamp 1607721120
transform 1 0 10948 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0774_
timestamp 1607721120
transform 1 0 9844 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_123
timestamp 1607721120
transform 1 0 12420 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1607721120
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1273_
timestamp 1607721120
transform 1 0 12512 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_15_143
timestamp 1607721120
transform 1 0 14260 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1274_
timestamp 1607721120
transform 1 0 14996 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1607721120
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_170
timestamp 1607721120
transform 1 0 16744 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_204
timestamp 1607721120
transform 1 0 19872 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_184
timestamp 1607721120
transform 1 0 18032 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_wb_clk_i
timestamp 1607721120
transform 1 0 18768 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1607721120
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1238_
timestamp 1607721120
transform 1 0 19044 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_215
timestamp 1607721120
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_wb_clk_i
timestamp 1607721120
transform 1 0 20608 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1318_
timestamp 1607721120
transform 1 0 21068 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1607721120
transform 1 0 24012 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_236
timestamp 1607721120
transform 1 0 22816 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1607721120
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1189_
timestamp 1607721120
transform 1 0 23644 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1607721120
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_261
timestamp 1607721120
transform 1 0 25116 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0857_
timestamp 1607721120
transform 1 0 25208 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_15_296
timestamp 1607721120
transform 1 0 28336 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1316_
timestamp 1607721120
transform 1 0 26588 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_15_313
timestamp 1607721120
transform 1 0 29900 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_304
timestamp 1607721120
transform 1 0 29072 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1607721120
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0880_
timestamp 1607721120
transform 1 0 29256 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_15_338
timestamp 1607721120
transform 1 0 32200 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_333
timestamp 1607721120
transform 1 0 31740 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_325
timestamp 1607721120
transform 1 0 31004 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0993_
timestamp 1607721120
transform 1 0 30636 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0923_
timestamp 1607721120
transform 1 0 31832 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_358
timestamp 1607721120
transform 1 0 34040 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _1140_
timestamp 1607721120
transform 1 0 32936 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_386
timestamp 1607721120
transform 1 0 36616 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1607721120
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1267_
timestamp 1607721120
transform 1 0 34868 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_15_402
timestamp 1607721120
transform 1 0 38088 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_398
timestamp 1607721120
transform 1 0 37720 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1130_
timestamp 1607721120
transform 1 0 38180 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_428
timestamp 1607721120
transform 1 0 40480 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_415
timestamp 1607721120
transform 1 0 39284 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1607721120
transform 1 0 40388 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_440
timestamp 1607721120
transform 1 0 41584 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1271_
timestamp 1607721120
transform 1 0 42136 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_15_465
timestamp 1607721120
transform 1 0 43884 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1191_
timestamp 1607721120
transform 1 0 44620 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_15_501
timestamp 1607721120
transform 1 0 47196 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_480
timestamp 1607721120
transform 1 0 45264 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1607721120
transform 1 0 46000 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1162_
timestamp 1607721120
transform 1 0 46092 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1263_
timestamp 1607721120
transform 1 0 48300 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_15_548
timestamp 1607721120
transform 1 0 51520 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_544
timestamp 1607721120
transform 1 0 51152 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_532
timestamp 1607721120
transform 1 0 50048 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_570
timestamp 1607721120
transform 1 0 53544 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_561
timestamp 1607721120
transform 1 0 52716 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_553
timestamp 1607721120
transform 1 0 51980 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1607721120
transform 1 0 51612 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1607721120
transform 1 0 51704 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0669_
timestamp 1607721120
transform 1 0 52900 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_15_582
timestamp 1607721120
transform 1 0 54648 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _1148_
timestamp 1607721120
transform 1 0 55384 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0728_
timestamp 1607721120
transform 1 0 54280 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_602
timestamp 1607721120
transform 1 0 56488 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1607721120
transform 1 0 57224 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1259_
timestamp 1607721120
transform 1 0 57316 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_15_630
timestamp 1607721120
transform 1 0 59064 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_660
timestamp 1607721120
transform 1 0 61824 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_654
timestamp 1607721120
transform 1 0 61272 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_642
timestamp 1607721120
transform 1 0 60168 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1607721120
transform -1 0 62192 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_15
timestamp 1607721120
transform 1 0 2484 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1607721120
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1607721120
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1231_
timestamp 1607721120
transform 1 0 2576 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1607721120
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1607721120
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1607721120
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1256_
timestamp 1607721120
transform 1 0 4416 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_16_55
timestamp 1607721120
transform 1 0 6164 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1234_
timestamp 1607721120
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1607721120
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1607721120
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_75
timestamp 1607721120
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_112
timestamp 1607721120
transform 1 0 11408 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1607721120
transform 1 0 10028 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1607721120
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0792_
timestamp 1607721120
transform 1 0 10764 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0769_
timestamp 1607721120
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1275_
timestamp 1607721120
transform 1 0 12144 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1607721120
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_139
timestamp 1607721120
transform 1 0 13892 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1607721120
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1125_
timestamp 1607721120
transform 1 0 15272 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_16_173
timestamp 1607721120
transform 1 0 17020 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_161
timestamp 1607721120
transform 1 0 15916 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1237_
timestamp 1607721120
transform 1 0 17296 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_16_205
timestamp 1607721120
transform 1 0 19964 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_183
timestamp 1607721120
transform 1 0 17940 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1242_
timestamp 1607721120
transform 1 0 18676 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_16_222
timestamp 1607721120
transform 1 0 21528 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1607721120
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1607721120
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0874_
timestamp 1607721120
transform 1 0 20884 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_16_243
timestamp 1607721120
transform 1 0 23460 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _0875_
timestamp 1607721120
transform 1 0 22264 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _0855_
timestamp 1607721120
transform 1 0 24196 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_267
timestamp 1607721120
transform 1 0 25668 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_255
timestamp 1607721120
transform 1 0 24564 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0856_
timestamp 1607721120
transform 1 0 25300 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_286
timestamp 1607721120
transform 1 0 27416 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1607721120
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1607721120
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0881_
timestamp 1607721120
transform 1 0 26588 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0877_
timestamp 1607721120
transform 1 0 28152 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_16_316
timestamp 1607721120
transform 1 0 30176 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_301
timestamp 1607721120
transform 1 0 28796 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1209_
timestamp 1607721120
transform 1 0 29532 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_16_341
timestamp 1607721120
transform 1 0 32476 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_328
timestamp 1607721120
transform 1 0 31280 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1607721120
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1106_
timestamp 1607721120
transform 1 0 30912 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0796_
timestamp 1607721120
transform 1 0 32108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1266_
timestamp 1607721120
transform 1 0 33212 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_16_376
timestamp 1607721120
transform 1 0 35696 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_368
timestamp 1607721120
transform 1 0 34960 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _1138_
timestamp 1607721120
transform 1 0 35788 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_402
timestamp 1607721120
transform 1 0 38088 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_389
timestamp 1607721120
transform 1 0 36892 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1607721120
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1128_
timestamp 1607721120
transform 1 0 37720 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_433
timestamp 1607721120
transform 1 0 40940 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1269_
timestamp 1607721120
transform 1 0 39192 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_16_450
timestamp 1607721120
transform 1 0 42504 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_441
timestamp 1607721120
transform 1 0 41676 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1199_
timestamp 1607721120
transform 1 0 41860 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_16_469
timestamp 1607721120
transform 1 0 44252 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_459
timestamp 1607721120
transform 1 0 43332 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1607721120
transform 1 0 43240 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1257_
timestamp 1607721120
transform 1 0 44988 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _0702_
timestamp 1607721120
transform 1 0 43608 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_16_496
timestamp 1607721120
transform 1 0 46736 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_511
timestamp 1607721120
transform 1 0 48116 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1607721120
transform 1 0 48852 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1261_
timestamp 1607721120
transform 1 0 48944 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1246_
timestamp 1607721120
transform 1 0 47472 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_16_547
timestamp 1607721120
transform 1 0 51428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_539
timestamp 1607721120
transform 1 0 50692 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_569
timestamp 1607721120
transform 1 0 53452 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1262_
timestamp 1607721120
transform 1 0 51704 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_16_588
timestamp 1607721120
transform 1 0 55200 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_577
timestamp 1607721120
transform 1 0 54188 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1607721120
transform 1 0 54464 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0673_
timestamp 1607721120
transform 1 0 54556 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_16_600
timestamp 1607721120
transform 1 0 56304 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1258_
timestamp 1607721120
transform 1 0 56396 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_16_632
timestamp 1607721120
transform 1 0 59248 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_620
timestamp 1607721120
transform 1 0 58144 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1146_
timestamp 1607721120
transform 1 0 58880 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_660
timestamp 1607721120
transform 1 0 61824 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_654
timestamp 1607721120
transform 1 0 61272 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_642
timestamp 1607721120
transform 1 0 60168 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_640
timestamp 1607721120
transform 1 0 59984 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1607721120
transform 1 0 60076 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1607721120
transform -1 0 62192 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_15
timestamp 1607721120
transform 1 0 2484 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1607721120
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1607721120
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0805_
timestamp 1607721120
transform 1 0 3036 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_17_28
timestamp 1607721120
transform 1 0 3680 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_4  _1235_
timestamp 1607721120
transform 1 0 4416 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_17_53
timestamp 1607721120
transform 1 0 5980 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1607721120
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0806_
timestamp 1607721120
transform 1 0 6808 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_17_91
timestamp 1607721120
transform 1 0 9476 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_76
timestamp 1607721120
transform 1 0 8096 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1232_
timestamp 1607721120
transform 1 0 8832 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_17_114
timestamp 1607721120
transform 1 0 11592 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 1607721120
transform 1 0 10580 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _0775_
timestamp 1607721120
transform 1 0 10948 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_17_137
timestamp 1607721120
transform 1 0 13708 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1607721120
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0793_
timestamp 1607721120
transform 1 0 12420 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_17_157
timestamp 1607721120
transform 1 0 15548 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _1126_
timestamp 1607721120
transform 1 0 14444 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_175
timestamp 1607721120
transform 1 0 17204 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_wb_clk_i
timestamp 1607721120
transform 1 0 16284 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1239_
timestamp 1607721120
transform 1 0 16560 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_17_197
timestamp 1607721120
transform 1 0 19228 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_184
timestamp 1607721120
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1607721120
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _1241_
timestamp 1607721120
transform 1 0 18400 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1229_
timestamp 1607721120
transform 1 0 19964 0 1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_17_219
timestamp 1607721120
transform 1 0 21252 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1221_
timestamp 1607721120
transform 1 0 21988 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_17_249
timestamp 1607721120
transform 1 0 24012 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_242
timestamp 1607721120
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_234
timestamp 1607721120
transform 1 0 22632 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1607721120
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0876_
timestamp 1607721120
transform 1 0 23644 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_272
timestamp 1607721120
transform 1 0 26128 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_261
timestamp 1607721120
transform 1 0 25116 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0870_
timestamp 1607721120
transform 1 0 24748 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1607721120
transform 1 0 25852 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_4  _1216_
timestamp 1607721120
transform 1 0 26864 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_17_306
timestamp 1607721120
transform 1 0 29256 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_297
timestamp 1607721120
transform 1 0 28428 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1607721120
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1207_
timestamp 1607721120
transform 1 0 29992 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_17_329
timestamp 1607721120
transform 1 0 31372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_321
timestamp 1607721120
transform 1 0 30636 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1214_
timestamp 1607721120
transform 1 0 31556 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_358
timestamp 1607721120
transform 1 0 34040 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_343
timestamp 1607721120
transform 1 0 32660 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1196_
timestamp 1607721120
transform 1 0 33396 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_17_382
timestamp 1607721120
transform 1 0 36248 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_374
timestamp 1607721120
transform 1 0 35512 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1607721120
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1268_
timestamp 1607721120
transform 1 0 36340 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _1194_
timestamp 1607721120
transform 1 0 34868 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_17_402
timestamp 1607721120
transform 1 0 38088 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_428
timestamp 1607721120
transform 1 0 40480 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_426
timestamp 1607721120
transform 1 0 40296 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_414
timestamp 1607721120
transform 1 0 39192 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1607721120
transform 1 0 40388 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1270_
timestamp 1607721120
transform 1 0 41584 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_17_479
timestamp 1607721120
transform 1 0 45172 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_459
timestamp 1607721120
transform 1 0 43332 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1200_
timestamp 1607721120
transform 1 0 44068 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_496
timestamp 1607721120
transform 1 0 46736 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_487
timestamp 1607721120
transform 1 0 45908 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1607721120
transform 1 0 46000 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0697_
timestamp 1607721120
transform 1 0 46092 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_17_525
timestamp 1607721120
transform 1 0 49404 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_512
timestamp 1607721120
transform 1 0 48208 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_508
timestamp 1607721120
transform 1 0 47840 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1154_
timestamp 1607721120
transform 1 0 48300 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_541
timestamp 1607721120
transform 1 0 50876 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0660_
timestamp 1607721120
transform 1 0 50508 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_570
timestamp 1607721120
transform 1 0 53544 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_562
timestamp 1607721120
transform 1 0 52808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1607721120
transform 1 0 51612 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1152_
timestamp 1607721120
transform 1 0 51704 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_587
timestamp 1607721120
transform 1 0 55108 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_579
timestamp 1607721120
transform 1 0 54372 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _1160_
timestamp 1607721120
transform 1 0 55384 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0661_
timestamp 1607721120
transform 1 0 53728 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_17_611
timestamp 1607721120
transform 1 0 57316 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_602
timestamp 1607721120
transform 1 0 56488 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1607721120
transform 1 0 57224 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1264_
timestamp 1607721120
transform 1 0 57684 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_17_634
timestamp 1607721120
transform 1 0 59432 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_658
timestamp 1607721120
transform 1 0 61640 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_646
timestamp 1607721120
transform 1 0 60536 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1607721120
transform -1 0 62192 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1607721120
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1607721120
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1607721120
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_44
timestamp 1607721120
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1607721120
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1607721120
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1607721120
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_60
timestamp 1607721120
transform 1 0 6624 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0802_
timestamp 1607721120
transform 1 0 5336 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _0779_
timestamp 1607721120
transform 1 0 7360 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1607721120
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1607721120
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_75
timestamp 1607721120
transform 1 0 8004 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_98
timestamp 1607721120
transform 1 0 10120 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1607721120
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1607721120
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0776_
timestamp 1607721120
transform 1 0 10856 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _0762_
timestamp 1607721120
transform 1 0 9752 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_135
timestamp 1607721120
transform 1 0 13524 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_120
timestamp 1607721120
transform 1 0 12144 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _0770_
timestamp 1607721120
transform 1 0 12880 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_18_154
timestamp 1607721120
transform 1 0 15272 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_147
timestamp 1607721120
transform 1 0 14628 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1607721120
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_169
timestamp 1607721120
transform 1 0 16652 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1224_
timestamp 1607721120
transform 1 0 16008 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1218_
timestamp 1607721120
transform 1 0 17388 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_18_192
timestamp 1607721120
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_184
timestamp 1607721120
transform 1 0 18032 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1219_
timestamp 1607721120
transform 1 0 18952 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_227
timestamp 1607721120
transform 1 0 21988 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_206
timestamp 1607721120
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1607721120
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1225_
timestamp 1607721120
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_242
timestamp 1607721120
transform 1 0 23368 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1227_
timestamp 1607721120
transform 1 0 22724 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1110_
timestamp 1607721120
transform 1 0 24104 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_267
timestamp 1607721120
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_262
timestamp 1607721120
transform 1 0 25208 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_254
timestamp 1607721120
transform 1 0 24472 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0878_
timestamp 1607721120
transform 1 0 25300 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_285
timestamp 1607721120
transform 1 0 27324 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_276
timestamp 1607721120
transform 1 0 26496 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1607721120
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _1215_
timestamp 1607721120
transform 1 0 28060 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__or2_4  _1212_
timestamp 1607721120
transform 1 0 26680 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_18_310
timestamp 1607721120
transform 1 0 29624 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _1208_
timestamp 1607721120
transform 1 0 30360 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_335
timestamp 1607721120
transform 1 0 31924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_327
timestamp 1607721120
transform 1 0 31188 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1607721120
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1204_
timestamp 1607721120
transform 1 0 32108 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_18_351
timestamp 1607721120
transform 1 0 33396 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1197_
timestamp 1607721120
transform 1 0 34132 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_387
timestamp 1607721120
transform 1 0 36708 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_368
timestamp 1607721120
transform 1 0 34960 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0729_
timestamp 1607721120
transform 1 0 36064 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_18_406
timestamp 1607721120
transform 1 0 38456 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_398
timestamp 1607721120
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_395
timestamp 1607721120
transform 1 0 37444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1607721120
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1272_
timestamp 1607721120
transform 1 0 38732 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_18_428
timestamp 1607721120
transform 1 0 40480 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_456
timestamp 1607721120
transform 1 0 43056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_448
timestamp 1607721120
transform 1 0 42320 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _1134_
timestamp 1607721120
transform 1 0 41216 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_471
timestamp 1607721120
transform 1 0 44436 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_463
timestamp 1607721120
transform 1 0 43700 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1607721120
transform 1 0 43240 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0698_
timestamp 1607721120
transform 1 0 44528 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _0688_
timestamp 1607721120
transform 1 0 43332 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1607721120
transform 1 0 47196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_486
timestamp 1607721120
transform 1 0 45816 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _0689_
timestamp 1607721120
transform 1 0 46552 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_18_520
timestamp 1607721120
transform 1 0 48944 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_513
timestamp 1607721120
transform 1 0 48300 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1607721120
transform 1 0 48852 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_548
timestamp 1607721120
transform 1 0 51520 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_533
timestamp 1607721120
transform 1 0 50140 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_528
timestamp 1607721120
transform 1 0 49680 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0655_
timestamp 1607721120
transform 1 0 49772 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _0651_
timestamp 1607721120
transform 1 0 50876 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_18_556
timestamp 1607721120
transform 1 0 52256 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0674_
timestamp 1607721120
transform 1 0 52440 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_18_572
timestamp 1607721120
transform 1 0 53728 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1607721120
transform 1 0 54464 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0656_
timestamp 1607721120
transform 1 0 54556 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_18_607
timestamp 1607721120
transform 1 0 56948 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_595
timestamp 1607721120
transform 1 0 55844 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _1156_
timestamp 1607721120
transform 1 0 57684 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_639
timestamp 1607721120
transform 1 0 59892 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_627
timestamp 1607721120
transform 1 0 58788 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_660
timestamp 1607721120
transform 1 0 61824 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_654
timestamp 1607721120
transform 1 0 61272 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_642
timestamp 1607721120
transform 1 0 60168 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1607721120
transform 1 0 60076 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1607721120
transform -1 0 62192 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1607721120
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1607721120
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1607721120
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1607721120
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1607721120
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1607721120
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1607721120
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1607721120
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1607721120
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1607721120
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0812_
timestamp 1607721120
transform 1 0 5152 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0811_
timestamp 1607721120
transform 1 0 4692 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1607721120
transform 1 0 7084 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1607721120
transform 1 0 5980 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_53
timestamp 1607721120
transform 1 0 5980 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1607721120
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0783_
timestamp 1607721120
transform 1 0 6808 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_20_89
timestamp 1607721120
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_77
timestamp 1607721120
transform 1 0 8188 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_87
timestamp 1607721120
transform 1 0 9108 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_81
timestamp 1607721120
transform 1 0 8556 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1607721120
transform 1 0 7452 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0763_
timestamp 1607721120
transform 1 0 9200 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1607721120
transform 1 0 11224 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_102
timestamp 1607721120
transform 1 0 10488 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_114
timestamp 1607721120
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_92
timestamp 1607721120
transform 1 0 9568 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1607721120
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0780_
timestamp 1607721120
transform 1 0 10304 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _0771_
timestamp 1607721120
transform 1 0 11408 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _0620_
timestamp 1607721120
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_126
timestamp 1607721120
transform 1 0 12696 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_137
timestamp 1607721120
transform 1 0 13708 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1607721120
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0765_
timestamp 1607721120
transform 1 0 12420 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _0764_
timestamp 1607721120
transform 1 0 13432 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_20_158
timestamp 1607721120
transform 1 0 15640 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1607721120
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_149
timestamp 1607721120
transform 1 0 14812 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_wb_clk_i
timestamp 1607721120
transform 1 0 15548 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1607721120
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0790_
timestamp 1607721120
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0742_
timestamp 1607721120
transform 1 0 14444 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_170
timestamp 1607721120
transform 1 0 16744 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_175
timestamp 1607721120
transform 1 0 17204 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1607721120
transform 1 0 15824 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1240_
timestamp 1607721120
transform 1 0 16560 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _1120_
timestamp 1607721120
transform 1 0 17112 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_186
timestamp 1607721120
transform 1 0 18216 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_195
timestamp 1607721120
transform 1 0 19044 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1607721120
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1607721120
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1230_
timestamp 1607721120
transform 1 0 18216 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1223_
timestamp 1607721120
transform 1 0 19780 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_4  _1114_
timestamp 1607721120
transform 1 0 18952 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_227
timestamp 1607721120
transform 1 0 21988 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_206
timestamp 1607721120
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_217
timestamp 1607721120
transform 1 0 21068 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1607721120
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1222_
timestamp 1607721120
transform 1 0 21804 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _1118_
timestamp 1607721120
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_242
timestamp 1607721120
transform 1 0 23368 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1607721120
transform 1 0 24012 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_242
timestamp 1607721120
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_234
timestamp 1607721120
transform 1 0 22632 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1607721120
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1195_
timestamp 1607721120
transform 1 0 24104 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0879_
timestamp 1607721120
transform 1 0 23644 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _0752_
timestamp 1607721120
transform 1 0 22724 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_20_267
timestamp 1607721120
transform 1 0 25668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_262
timestamp 1607721120
transform 1 0 25208 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_254
timestamp 1607721120
transform 1 0 24472 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_265
timestamp 1607721120
transform 1 0 25484 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_261
timestamp 1607721120
transform 1 0 25116 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1193_
timestamp 1607721120
transform 1 0 25300 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1116_
timestamp 1607721120
transform 1 0 25576 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_288
timestamp 1607721120
transform 1 0 27600 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1607721120
transform 1 0 28060 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_278
timestamp 1607721120
transform 1 0 26680 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1607721120
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1217_
timestamp 1607721120
transform 1 0 26496 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1211_
timestamp 1607721120
transform 1 0 28336 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _1210_
timestamp 1607721120
transform 1 0 27416 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_20_311
timestamp 1607721120
transform 1 0 29716 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_303
timestamp 1607721120
transform 1 0 28980 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_312
timestamp 1607721120
transform 1 0 29808 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_306
timestamp 1607721120
transform 1 0 29256 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1607721120
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _1112_
timestamp 1607721120
transform 1 0 29900 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0644_
timestamp 1607721120
transform 1 0 29440 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_333
timestamp 1607721120
transform 1 0 31740 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_325
timestamp 1607721120
transform 1 0 31004 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_327
timestamp 1607721120
transform 1 0 31188 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1607721120
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1213_
timestamp 1607721120
transform 1 0 30544 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _1205_
timestamp 1607721120
transform 1 0 32108 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _1198_
timestamp 1607721120
transform 1 0 31924 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_20_363
timestamp 1607721120
transform 1 0 34500 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_346
timestamp 1607721120
transform 1 0 32936 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_365
timestamp 1607721120
transform 1 0 34684 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_361
timestamp 1607721120
transform 1 0 34316 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1607721120
transform 1 0 33212 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _1203_
timestamp 1607721120
transform 1 0 33672 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_19_372
timestamp 1607721120
transform 1 0 35328 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_367
timestamp 1607721120
transform 1 0 34868 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1607721120
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0714_
timestamp 1607721120
transform 1 0 34960 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_379
timestamp 1607721120
transform 1 0 35972 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_375
timestamp 1607721120
transform 1 0 35604 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _0724_
timestamp 1607721120
transform 1 0 36064 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0719_
timestamp 1607721120
transform 1 0 36064 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_20_387
timestamp 1607721120
transform 1 0 36708 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_387
timestamp 1607721120
transform 1 0 36708 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_395
timestamp 1607721120
transform 1 0 37444 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_402
timestamp 1607721120
transform 1 0 38088 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1607721120
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0720_
timestamp 1607721120
transform 1 0 37720 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_4  _0715_
timestamp 1607721120
transform 1 0 37444 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_20_424
timestamp 1607721120
transform 1 0 40112 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_412
timestamp 1607721120
transform 1 0 39008 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_426
timestamp 1607721120
transform 1 0 40296 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_414
timestamp 1607721120
transform 1 0 39192 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1607721120
transform 1 0 40388 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0710_
timestamp 1607721120
transform 1 0 40480 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_20_446
timestamp 1607721120
transform 1 0 42136 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_436
timestamp 1607721120
transform 1 0 41216 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_451
timestamp 1607721120
transform 1 0 42596 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_443
timestamp 1607721120
transform 1 0 41860 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_435
timestamp 1607721120
transform 1 0 41124 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_wb_clk_i
timestamp 1607721120
transform 1 0 42872 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1206_
timestamp 1607721120
transform 1 0 41492 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0693_
timestamp 1607721120
transform 1 0 41952 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_20_471
timestamp 1607721120
transform 1 0 44436 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_459
timestamp 1607721120
transform 1 0 43332 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_457
timestamp 1607721120
transform 1 0 43148 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_471
timestamp 1607721120
transform 1 0 44436 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_wb_clk_i
timestamp 1607721120
transform 1 0 45172 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1607721120
transform 1 0 43240 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _1192_
timestamp 1607721120
transform 1 0 43332 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _0694_
timestamp 1607721120
transform 1 0 44528 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_20_486
timestamp 1607721120
transform 1 0 45816 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_482
timestamp 1607721120
transform 1 0 45448 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_wb_clk_i
timestamp 1607721120
transform 1 0 46552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1607721120
transform 1 0 46000 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1247_
timestamp 1607721120
transform 1 0 46092 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _0690_
timestamp 1607721120
transform 1 0 46828 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_20_511
timestamp 1607721120
transform 1 0 48116 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_515
timestamp 1607721120
transform 1 0 48484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_503
timestamp 1607721120
transform 1 0 47380 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1607721120
transform 1 0 48852 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0684_
timestamp 1607721120
transform 1 0 48944 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _0654_
timestamp 1607721120
transform 1 0 48116 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_542
timestamp 1607721120
transform 1 0 50968 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_534
timestamp 1607721120
transform 1 0 50232 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_541
timestamp 1607721120
transform 1 0 50876 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_533
timestamp 1607721120
transform 1 0 50140 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_527
timestamp 1607721120
transform 1 0 49588 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _0683_
timestamp 1607721120
transform 1 0 50232 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0665_
timestamp 1607721120
transform 1 0 51060 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_20_550
timestamp 1607721120
transform 1 0 51704 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_558
timestamp 1607721120
transform 1 0 52440 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_550
timestamp 1607721120
transform 1 0 51704 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1607721120
transform 1 0 51612 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0670_
timestamp 1607721120
transform 1 0 52440 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _0666_
timestamp 1607721120
transform 1 0 52624 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1607721120
transform 1 0 55292 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_581
timestamp 1607721120
transform 1 0 54556 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_572
timestamp 1607721120
transform 1 0 53728 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_574
timestamp 1607721120
transform 1 0 53912 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1607721120
transform 1 0 54464 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0664_
timestamp 1607721120
transform 1 0 54648 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0662_
timestamp 1607721120
transform 1 0 54648 0 1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_20_613
timestamp 1607721120
transform 1 0 57500 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1607721120
transform 1 0 56396 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_611
timestamp 1607721120
transform 1 0 57316 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_608
timestamp 1607721120
transform 1 0 57040 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_596
timestamp 1607721120
transform 1 0 55936 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1607721120
transform 1 0 57224 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_637
timestamp 1607721120
transform 1 0 59708 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_625
timestamp 1607721120
transform 1 0 58604 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_619
timestamp 1607721120
transform 1 0 58052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1260_
timestamp 1607721120
transform 1 0 58328 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_20_660
timestamp 1607721120
transform 1 0 61824 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_654
timestamp 1607721120
transform 1 0 61272 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_642
timestamp 1607721120
transform 1 0 60168 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_653
timestamp 1607721120
transform 1 0 61180 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_641
timestamp 1607721120
transform 1 0 60076 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1607721120
transform 1 0 60076 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1607721120
transform -1 0 62192 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1607721120
transform -1 0 62192 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1607721120
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1607721120
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1607721120
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_43
timestamp 1607721120
transform 1 0 5060 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_39
timestamp 1607721120
transform 1 0 4692 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1607721120
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _0807_
timestamp 1607721120
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_53
timestamp 1607721120
transform 1 0 5980 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1607721120
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0803_
timestamp 1607721120
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_83
timestamp 1607721120
transform 1 0 8740 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_71
timestamp 1607721120
transform 1 0 7636 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1607721120
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_99
timestamp 1607721120
transform 1 0 10212 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_95
timestamp 1607721120
transform 1 0 9844 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _0784_
timestamp 1607721120
transform 1 0 10304 0 1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_21_132
timestamp 1607721120
transform 1 0 13248 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1607721120
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0794_
timestamp 1607721120
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1607721120
transform 1 0 14812 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _0799_
timestamp 1607721120
transform 1 0 13984 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1607721120
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_173
timestamp 1607721120
transform 1 0 17020 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_161
timestamp 1607721120
transform 1 0 15916 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_192
timestamp 1607721120
transform 1 0 18768 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_184
timestamp 1607721120
transform 1 0 18032 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1607721120
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1277_
timestamp 1607721120
transform 1 0 19504 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _1243_
timestamp 1607721120
transform 1 0 18124 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_21_219
timestamp 1607721120
transform 1 0 21252 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1228_
timestamp 1607721120
transform 1 0 21988 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_251
timestamp 1607721120
transform 1 0 24196 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_245
timestamp 1607721120
transform 1 0 23644 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_236
timestamp 1607721120
transform 1 0 22816 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1607721120
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_267
timestamp 1607721120
transform 1 0 25668 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_259
timestamp 1607721120
transform 1 0 24932 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1278_
timestamp 1607721120
transform 1 0 25852 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__and2_4  _0748_
timestamp 1607721120
transform 1 0 24288 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_21_288
timestamp 1607721120
transform 1 0 27600 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_314
timestamp 1607721120
transform 1 0 29992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_306
timestamp 1607721120
transform 1 0 29256 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_304
timestamp 1607721120
transform 1 0 29072 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_300
timestamp 1607721120
transform 1 0 28704 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1607721120
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1280_
timestamp 1607721120
transform 1 0 30176 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_21_335
timestamp 1607721120
transform 1 0 31924 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_362
timestamp 1607721120
transform 1 0 34408 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_350
timestamp 1607721120
transform 1 0 33304 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0737_
timestamp 1607721120
transform 1 0 32660 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_21_379
timestamp 1607721120
transform 1 0 35972 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_371
timestamp 1607721120
transform 1 0 35236 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1607721120
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0725_
timestamp 1607721120
transform 1 0 36156 0 1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _0621_
timestamp 1607721120
transform 1 0 34868 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_395
timestamp 1607721120
transform 1 0 37444 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0716_
timestamp 1607721120
transform 1 0 38180 0 1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_21_428
timestamp 1607721120
transform 1 0 40480 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_425
timestamp 1607721120
transform 1 0 40204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_417
timestamp 1607721120
transform 1 0 39468 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1607721120
transform 1 0 40388 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_452
timestamp 1607721120
transform 1 0 42688 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_440
timestamp 1607721120
transform 1 0 41584 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_464
timestamp 1607721120
transform 1 0 43792 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0703_
timestamp 1607721120
transform 1 0 43976 0 1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_21_498
timestamp 1607721120
transform 1 0 46920 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_480
timestamp 1607721120
transform 1 0 45264 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1607721120
transform 1 0 46000 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1248_
timestamp 1607721120
transform 1 0 46092 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_524
timestamp 1607721120
transform 1 0 49312 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_512
timestamp 1607721120
transform 1 0 48208 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_506
timestamp 1607721120
transform 1 0 47656 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0682_
timestamp 1607721120
transform 1 0 47840 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0681_
timestamp 1607721120
transform 1 0 48944 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_541
timestamp 1607721120
transform 1 0 50876 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_536
timestamp 1607721120
transform 1 0 50416 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0645_
timestamp 1607721120
transform 1 0 50508 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_559
timestamp 1607721120
transform 1 0 52532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1607721120
transform 1 0 51612 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0675_
timestamp 1607721120
transform 1 0 51704 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_581
timestamp 1607721120
transform 1 0 54556 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_571
timestamp 1607721120
transform 1 0 53636 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0667_
timestamp 1607721120
transform 1 0 53728 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _0657_
timestamp 1607721120
transform 1 0 55292 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_21_611
timestamp 1607721120
transform 1 0 57316 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_598
timestamp 1607721120
transform 1 0 56120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1607721120
transform 1 0 57224 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_635
timestamp 1607721120
transform 1 0 59524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_623
timestamp 1607721120
transform 1 0 58420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_659
timestamp 1607721120
transform 1 0 61732 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_647
timestamp 1607721120
transform 1 0 60628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1607721120
transform -1 0 62192 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1607721120
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1607721120
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1607721120
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_32
timestamp 1607721120
transform 1 0 4048 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1607721120
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1607721120
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1326_
timestamp 1607721120
transform 1 0 4600 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_22_57
timestamp 1607721120
transform 1 0 6348 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1327_
timestamp 1607721120
transform 1 0 7084 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_22_84
timestamp 1607721120
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_107
timestamp 1607721120
transform 1 0 10948 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_99
timestamp 1607721120
transform 1 0 10212 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_93
timestamp 1607721120
transform 1 0 9660 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1607721120
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0795_
timestamp 1607721120
transform 1 0 10304 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_22_134
timestamp 1607721120
transform 1 0 13432 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1329_
timestamp 1607721120
transform 1 0 11684 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_22_158
timestamp 1607721120
transform 1 0 15640 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1607721120
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_146
timestamp 1607721120
transform 1 0 14536 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1607721120
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0787_
timestamp 1607721120
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_166
timestamp 1607721120
transform 1 0 16376 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1276_
timestamp 1607721120
transform 1 0 16652 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_22_196
timestamp 1607721120
transform 1 0 19136 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1607721120
transform 1 0 18400 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _0743_
timestamp 1607721120
transform 1 0 19412 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1607721120
transform 1 0 20884 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_206
timestamp 1607721120
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1607721120
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0744_
timestamp 1607721120
transform 1 0 21620 0 -1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_22_237
timestamp 1607721120
transform 1 0 22908 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0749_
timestamp 1607721120
transform 1 0 23644 0 -1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_22_271
timestamp 1607721120
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_259
timestamp 1607721120
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_285
timestamp 1607721120
transform 1 0 27324 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_276
timestamp 1607721120
transform 1 0 26496 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1607721120
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1226_
timestamp 1607721120
transform 1 0 26680 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_22_315
timestamp 1607721120
transform 1 0 30084 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_297
timestamp 1607721120
transform 1 0 28428 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _0738_
timestamp 1607721120
transform 1 0 28796 0 -1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_22_337
timestamp 1607721120
transform 1 0 32108 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_335
timestamp 1607721120
transform 1 0 31924 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_327
timestamp 1607721120
transform 1 0 31188 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1607721120
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0735_
timestamp 1607721120
transform 1 0 30820 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_353
timestamp 1607721120
transform 1 0 33580 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_345
timestamp 1607721120
transform 1 0 32844 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0813_
timestamp 1607721120
transform 1 0 32936 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _0731_
timestamp 1607721120
transform 1 0 34316 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_22_385
timestamp 1607721120
transform 1 0 36524 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_370
timestamp 1607721120
transform 1 0 35144 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1201_
timestamp 1607721120
transform 1 0 35880 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_22_404
timestamp 1607721120
transform 1 0 38272 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_398
timestamp 1607721120
transform 1 0 37720 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1607721120
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0708_
timestamp 1607721120
transform 1 0 37904 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_426
timestamp 1607721120
transform 1 0 40296 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _0711_
timestamp 1607721120
transform 1 0 39008 0 -1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_22_450
timestamp 1607721120
transform 1 0 42504 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_438
timestamp 1607721120
transform 1 0 41400 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_466
timestamp 1607721120
transform 1 0 43976 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_459
timestamp 1607721120
transform 1 0 43332 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1607721120
transform 1 0 43240 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1356_
timestamp 1607721120
transform 1 0 44712 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0677_
timestamp 1607721120
transform 1 0 43608 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_493
timestamp 1607721120
transform 1 0 46460 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0622_
timestamp 1607721120
transform 1 0 47196 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_520
timestamp 1607721120
transform 1 0 48944 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_517
timestamp 1607721120
transform 1 0 48668 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_505
timestamp 1607721120
transform 1 0 47564 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1607721120
transform 1 0 48852 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_532
timestamp 1607721120
transform 1 0 50048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1351_
timestamp 1607721120
transform 1 0 50232 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_22_570
timestamp 1607721120
transform 1 0 53544 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_553
timestamp 1607721120
transform 1 0 51980 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0671_
timestamp 1607721120
transform 1 0 52716 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_578
timestamp 1607721120
transform 1 0 54280 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1607721120
transform 1 0 54464 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1353_
timestamp 1607721120
transform 1 0 54556 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_22_600
timestamp 1607721120
transform 1 0 56304 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1355_
timestamp 1607721120
transform 1 0 57040 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_639
timestamp 1607721120
transform 1 0 59892 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_627
timestamp 1607721120
transform 1 0 58788 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_660
timestamp 1607721120
transform 1 0 61824 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_654
timestamp 1607721120
transform 1 0 61272 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_642
timestamp 1607721120
transform 1 0 60168 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1607721120
transform 1 0 60076 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1607721120
transform -1 0 62192 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1607721120
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1607721120
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1607721120
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_45
timestamp 1607721120
transform 1 0 5244 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_39
timestamp 1607721120
transform 1 0 4692 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1607721120
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1607721120
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_53
timestamp 1607721120
transform 1 0 5980 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1607721120
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1328_
timestamp 1607721120
transform 1 0 6992 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _0804_
timestamp 1607721120
transform 1 0 5336 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_23_83
timestamp 1607721120
transform 1 0 8740 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_114
timestamp 1607721120
transform 1 0 11592 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_95
timestamp 1607721120
transform 1 0 9844 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0788_
timestamp 1607721120
transform 1 0 10948 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1607721120
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1330_
timestamp 1607721120
transform 1 0 12420 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_23_157
timestamp 1607721120
transform 1 0 15548 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_150
timestamp 1607721120
transform 1 0 14904 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_142
timestamp 1607721120
transform 1 0 14168 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0759_
timestamp 1607721120
transform 1 0 15180 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1607721120
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_174
timestamp 1607721120
transform 1 0 17112 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0777_
timestamp 1607721120
transform 1 0 16284 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_188
timestamp 1607721120
transform 1 0 18400 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1607721120
transform 1 0 18032 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1607721120
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1279_
timestamp 1607721120
transform 1 0 18492 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_23_220
timestamp 1607721120
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1607721120
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _0757_
timestamp 1607721120
transform 1 0 21528 0 1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_23_236
timestamp 1607721120
transform 1 0 22816 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1607721120
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0758_
timestamp 1607721120
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1607721120
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_254
timestamp 1607721120
transform 1 0 24472 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0746_
timestamp 1607721120
transform 1 0 25208 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_23_294
timestamp 1607721120
transform 1 0 28152 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_282
timestamp 1607721120
transform 1 0 27048 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_277
timestamp 1607721120
transform 1 0 26588 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1607721120
transform 1 0 26772 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0732_
timestamp 1607721120
transform 1 0 27784 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_318
timestamp 1607721120
transform 1 0 30360 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_306
timestamp 1607721120
transform 1 0 29256 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_302
timestamp 1607721120
transform 1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1607721120
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_341
timestamp 1607721120
transform 1 0 32476 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_329
timestamp 1607721120
transform 1 0 31372 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1220_
timestamp 1607721120
transform 1 0 30728 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0705_
timestamp 1607721120
transform 1 0 32108 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_358
timestamp 1607721120
transform 1 0 34040 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0819_
timestamp 1607721120
transform 1 0 33212 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_387
timestamp 1607721120
transform 1 0 36708 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_379
timestamp 1607721120
transform 1 0 35972 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_367
timestamp 1607721120
transform 1 0 34868 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1607721120
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0730_
timestamp 1607721120
transform 1 0 36800 0 1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__and3_4  _0726_
timestamp 1607721120
transform 1 0 35144 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_402
timestamp 1607721120
transform 1 0 38088 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0709_
timestamp 1607721120
transform 1 0 38824 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_428
timestamp 1607721120
transform 1 0 40480 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_426
timestamp 1607721120
transform 1 0 40296 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_414
timestamp 1607721120
transform 1 0 39192 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1607721120
transform 1 0 40388 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_452
timestamp 1607721120
transform 1 0 42688 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_440
timestamp 1607721120
transform 1 0 41584 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_478
timestamp 1607721120
transform 1 0 45080 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_463
timestamp 1607721120
transform 1 0 43700 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_458
timestamp 1607721120
transform 1 0 43240 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0696_
timestamp 1607721120
transform 1 0 44436 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0676_
timestamp 1607721120
transform 1 0 43332 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_496
timestamp 1607721120
transform 1 0 46736 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_486
timestamp 1607721120
transform 1 0 45816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1607721120
transform 1 0 46000 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1245_
timestamp 1607721120
transform 1 0 46092 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_23_520
timestamp 1607721120
transform 1 0 48944 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_508
timestamp 1607721120
transform 1 0 47840 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0639_
timestamp 1607721120
transform 1 0 47472 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_548
timestamp 1607721120
transform 1 0 51520 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_544
timestamp 1607721120
transform 1 0 51152 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_532
timestamp 1607721120
transform 1 0 50048 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_569
timestamp 1607721120
transform 1 0 53452 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1607721120
transform 1 0 51612 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1352_
timestamp 1607721120
transform 1 0 51704 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_23_581
timestamp 1607721120
transform 1 0 54556 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _0663_
timestamp 1607721120
transform 1 0 54924 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_611
timestamp 1607721120
transform 1 0 57316 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_606
timestamp 1607721120
transform 1 0 56856 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_594
timestamp 1607721120
transform 1 0 55752 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1607721120
transform 1 0 57224 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_635
timestamp 1607721120
transform 1 0 59524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_623
timestamp 1607721120
transform 1 0 58420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_659
timestamp 1607721120
transform 1 0 61732 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_647
timestamp 1607721120
transform 1 0 60628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1607721120
transform -1 0 62192 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1607721120
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1607721120
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1607721120
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_44
timestamp 1607721120
transform 1 0 5152 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1607721120
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1607721120
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1607721120
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_67
timestamp 1607721120
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_55
timestamp 1607721120
transform 1 0 6164 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0808_
timestamp 1607721120
transform 1 0 5520 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1607721120
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_76
timestamp 1607721120
transform 1 0 8096 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0800_
timestamp 1607721120
transform 1 0 7452 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_24_110
timestamp 1607721120
transform 1 0 11224 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_105
timestamp 1607721120
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1607721120
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1607721120
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0786_
timestamp 1607721120
transform 1 0 10856 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_128
timestamp 1607721120
transform 1 0 12880 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_118
timestamp 1607721120
transform 1 0 11960 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0785_
timestamp 1607721120
transform 1 0 12052 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0782_
timestamp 1607721120
transform 1 0 13616 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1607721120
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1607721120
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_143
timestamp 1607721120
transform 1 0 14260 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1607721120
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0760_
timestamp 1607721120
transform 1 0 15456 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_160
timestamp 1607721120
transform 1 0 15824 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1335_
timestamp 1607721120
transform 1 0 16928 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_24_203
timestamp 1607721120
transform 1 0 19780 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_191
timestamp 1607721120
transform 1 0 18676 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1190_
timestamp 1607721120
transform 1 0 19412 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_227
timestamp 1607721120
transform 1 0 21988 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1607721120
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_211
timestamp 1607721120
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1607721120
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1607721120
transform 1 0 23460 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0753_
timestamp 1607721120
transform 1 0 22172 0 -1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__and3_4  _0750_
timestamp 1607721120
transform 1 0 24196 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_272
timestamp 1607721120
transform 1 0 26128 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_260
timestamp 1607721120
transform 1 0 25024 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_286
timestamp 1607721120
transform 1 0 27416 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_276
timestamp 1607721120
transform 1 0 26496 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1607721120
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0733_
timestamp 1607721120
transform 1 0 27048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_319
timestamp 1607721120
transform 1 0 30452 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_307
timestamp 1607721120
transform 1 0 29348 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _0739_
timestamp 1607721120
transform 1 0 28520 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_337
timestamp 1607721120
transform 1 0 32108 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_328
timestamp 1607721120
transform 1 0 31280 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_323
timestamp 1607721120
transform 1 0 30820 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1607721120
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0736_
timestamp 1607721120
transform 1 0 30912 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_364
timestamp 1607721120
transform 1 0 34592 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1325_
timestamp 1607721120
transform 1 0 32844 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_24_376
timestamp 1607721120
transform 1 0 35696 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__and3_4  _0721_
timestamp 1607721120
transform 1 0 36064 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_24_398
timestamp 1607721120
transform 1 0 37720 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_389
timestamp 1607721120
transform 1 0 36892 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1607721120
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0712_
timestamp 1607721120
transform 1 0 38272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_425
timestamp 1607721120
transform 1 0 40204 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_413
timestamp 1607721120
transform 1 0 39100 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_449
timestamp 1607721120
transform 1 0 42412 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_437
timestamp 1607721120
transform 1 0 41308 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_469
timestamp 1607721120
transform 1 0 44252 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_459
timestamp 1607721120
transform 1 0 43332 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_457
timestamp 1607721120
transform 1 0 43148 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1607721120
transform 1 0 43240 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0704_
timestamp 1607721120
transform 1 0 43424 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _0695_
timestamp 1607721120
transform 1 0 44988 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_498
timestamp 1607721120
transform 1 0 46920 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_486
timestamp 1607721120
transform 1 0 45816 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _0691_
timestamp 1607721120
transform 1 0 47288 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_511
timestamp 1607721120
transform 1 0 48116 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1607721120
transform 1 0 48852 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0685_
timestamp 1607721120
transform 1 0 48944 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_541
timestamp 1607721120
transform 1 0 50876 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_529
timestamp 1607721120
transform 1 0 49772 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0672_
timestamp 1607721120
transform 1 0 50968 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_24_564
timestamp 1607721120
transform 1 0 52992 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_549
timestamp 1607721120
transform 1 0 51612 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0668_
timestamp 1607721120
transform 1 0 52348 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_24_593
timestamp 1607721120
transform 1 0 55660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_581
timestamp 1607721120
transform 1 0 54556 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_576
timestamp 1607721120
transform 1 0 54096 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1607721120
transform 1 0 54464 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_614
timestamp 1607721120
transform 1 0 57592 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_602
timestamp 1607721120
transform 1 0 56488 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0640_
timestamp 1607721120
transform 1 0 55844 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_24_638
timestamp 1607721120
transform 1 0 59800 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_626
timestamp 1607721120
transform 1 0 58696 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_660
timestamp 1607721120
transform 1 0 61824 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_654
timestamp 1607721120
transform 1 0 61272 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_642
timestamp 1607721120
transform 1 0 60168 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1607721120
transform 1 0 60076 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1607721120
transform -1 0 62192 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1607721120
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1607721120
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1607721120
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1607721120
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1607721120
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1607721120
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1607721120
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1607721120
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1607721120
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1607721120
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1607721120
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1607721120
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1607721120
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_134
timestamp 1607721120
transform 1 0 13432 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1607721120
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1607721120
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0781_
timestamp 1607721120
transform 1 0 12604 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1607721120
transform 1 0 14812 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0778_
timestamp 1607721120
transform 1 0 14168 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1607721120
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_173
timestamp 1607721120
transform 1 0 17020 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_161
timestamp 1607721120
transform 1 0 15916 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _0766_
timestamp 1607721120
transform 1 0 16192 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_25_205
timestamp 1607721120
transform 1 0 19964 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1607721120
transform 1 0 18860 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1607721120
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0772_
timestamp 1607721120
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_219
timestamp 1607721120
transform 1 0 21252 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_211
timestamp 1607721120
transform 1 0 20516 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0756_
timestamp 1607721120
transform 1 0 20608 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _0754_
timestamp 1607721120
transform 1 0 21988 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_236
timestamp 1607721120
transform 1 0 22816 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1607721120
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1337_
timestamp 1607721120
transform 1 0 23644 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_25_264
timestamp 1607721120
transform 1 0 25392 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1607721120
transform 1 0 28060 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_276
timestamp 1607721120
transform 1 0 26496 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0745_
timestamp 1607721120
transform 1 0 27232 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1607721120
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1340_
timestamp 1607721120
transform 1 0 29256 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1607721120
transform 1 0 32108 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_325
timestamp 1607721120
transform 1 0 31004 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_358
timestamp 1607721120
transform 1 0 34040 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_353
timestamp 1607721120
transform 1 0 33580 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_349
timestamp 1607721120
transform 1 0 33212 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0706_
timestamp 1607721120
transform 1 0 33672 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_374
timestamp 1607721120
transform 1 0 35512 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1607721120
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1343_
timestamp 1607721120
transform 1 0 36248 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _0722_
timestamp 1607721120
transform 1 0 34868 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_25_401
timestamp 1607721120
transform 1 0 37996 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0717_
timestamp 1607721120
transform 1 0 38732 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_428
timestamp 1607721120
transform 1 0 40480 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_426
timestamp 1607721120
transform 1 0 40296 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_418
timestamp 1607721120
transform 1 0 39560 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1607721120
transform 1 0 40388 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_446
timestamp 1607721120
transform 1 0 42136 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_440
timestamp 1607721120
transform 1 0 41584 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0700_
timestamp 1607721120
transform 1 0 42872 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0678_
timestamp 1607721120
transform 1 0 41768 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_478
timestamp 1607721120
transform 1 0 45080 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_461
timestamp 1607721120
transform 1 0 43516 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0699_
timestamp 1607721120
transform 1 0 44252 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_496
timestamp 1607721120
transform 1 0 46736 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_486
timestamp 1607721120
transform 1 0 45816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1607721120
transform 1 0 46000 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0692_
timestamp 1607721120
transform 1 0 46092 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_25_508
timestamp 1607721120
transform 1 0 47840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1349_
timestamp 1607721120
transform 1 0 48024 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_25_541
timestamp 1607721120
transform 1 0 50876 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1607721120
transform 1 0 49772 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_562
timestamp 1607721120
transform 1 0 52808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_550
timestamp 1607721120
transform 1 0 51704 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1607721120
transform 1 0 51612 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_586
timestamp 1607721120
transform 1 0 55016 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_574
timestamp 1607721120
transform 1 0 53912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0658_
timestamp 1607721120
transform 1 0 55568 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_25_611
timestamp 1607721120
transform 1 0 57316 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_607
timestamp 1607721120
transform 1 0 56948 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_599
timestamp 1607721120
transform 1 0 56212 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1607721120
transform 1 0 57224 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_635
timestamp 1607721120
transform 1 0 59524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_623
timestamp 1607721120
transform 1 0 58420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_659
timestamp 1607721120
transform 1 0 61732 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_647
timestamp 1607721120
transform 1 0 60628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1607721120
transform -1 0 62192 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1607721120
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1607721120
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1607721120
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1607721120
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1607721120
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1607721120
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1607721120
transform 1 0 5152 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1607721120
transform 1 0 4048 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1607721120
transform 1 0 3588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1607721120
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1607721120
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1607721120
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1607721120
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1607721120
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_63
timestamp 1607721120
transform 1 0 6900 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_56
timestamp 1607721120
transform 1 0 6256 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1607721120
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1607721120
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1607721120
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_87
timestamp 1607721120
transform 1 0 9108 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_75
timestamp 1607721120
transform 1 0 8004 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1607721120
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_106
timestamp 1607721120
transform 1 0 10856 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_94
timestamp 1607721120
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_113
timestamp 1607721120
transform 1 0 11500 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_105
timestamp 1607721120
transform 1 0 10764 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1607721120
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1607721120
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1607721120
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 1607721120
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_118
timestamp 1607721120
transform 1 0 11960 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_135
timestamp 1607721120
transform 1 0 13524 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1607721120
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1332_
timestamp 1607721120
transform 1 0 12788 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1331_
timestamp 1607721120
transform 1 0 11776 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_27_156
timestamp 1607721120
transform 1 0 15456 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_154
timestamp 1607721120
transform 1 0 15272 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_146
timestamp 1607721120
transform 1 0 14536 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_147
timestamp 1607721120
transform 1 0 14628 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1607721120
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1607721120
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0773_
timestamp 1607721120
transform 1 0 15272 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_27_177
timestamp 1607721120
transform 1 0 17388 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_168
timestamp 1607721120
transform 1 0 16560 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_161
timestamp 1607721120
transform 1 0 15916 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1333_
timestamp 1607721120
transform 1 0 16652 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _0761_
timestamp 1607721120
transform 1 0 16744 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_27_185
timestamp 1607721120
transform 1 0 18124 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_203
timestamp 1607721120
transform 1 0 19780 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_188
timestamp 1607721120
transform 1 0 18400 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1607721120
transform 1 0 18216 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1334_
timestamp 1607721120
transform 1 0 18308 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _0767_
timestamp 1607721120
transform 1 0 19136 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_27_214
timestamp 1607721120
transform 1 0 20792 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_206
timestamp 1607721120
transform 1 0 20056 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1607721120
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_211
timestamp 1607721120
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1607721120
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_227
timestamp 1607721120
transform 1 0 21988 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1607721120
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1607721120
transform 1 0 21068 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0755_
timestamp 1607721120
transform 1 0 21344 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_27_218
timestamp 1607721120
transform 1 0 21160 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_240
timestamp 1607721120
transform 1 0 23184 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_230
timestamp 1607721120
transform 1 0 22264 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1607721120
transform 1 0 23920 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1338_
timestamp 1607721120
transform 1 0 24012 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1336_
timestamp 1607721120
transform 1 0 22724 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _0751_
timestamp 1607721120
transform 1 0 22540 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_27_268
timestamp 1607721120
transform 1 0 25760 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_274
timestamp 1607721120
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_266
timestamp 1607721120
transform 1 0 25576 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_254
timestamp 1607721120
transform 1 0 24472 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_288
timestamp 1607721120
transform 1 0 27600 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_280
timestamp 1607721120
transform 1 0 26864 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_276
timestamp 1607721120
transform 1 0 26496 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_288
timestamp 1607721120
transform 1 0 27600 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1607721120
transform 1 0 26496 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1607721120
transform 1 0 26772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1607721120
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1339_
timestamp 1607721120
transform 1 0 27692 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _0740_
timestamp 1607721120
transform 1 0 27876 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_27_311
timestamp 1607721120
transform 1 0 29716 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_298
timestamp 1607721120
transform 1 0 28520 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_308
timestamp 1607721120
transform 1 0 29440 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1607721120
transform 1 0 29624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0734_
timestamp 1607721120
transform 1 0 30176 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_27_342
timestamp 1607721120
transform 1 0 32568 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_335
timestamp 1607721120
transform 1 0 31924 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_323
timestamp 1607721120
transform 1 0 30820 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_337
timestamp 1607721120
transform 1 0 32108 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_335
timestamp 1607721120
transform 1 0 31924 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_323
timestamp 1607721120
transform 1 0 30820 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1607721120
transform 1 0 32476 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1607721120
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1341_
timestamp 1607721120
transform 1 0 32384 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_27_364
timestamp 1607721120
transform 1 0 34592 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_354
timestamp 1607721120
transform 1 0 33672 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_359
timestamp 1607721120
transform 1 0 34132 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0727_
timestamp 1607721120
transform 1 0 33948 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_27_380
timestamp 1607721120
transform 1 0 36064 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_386
timestamp 1607721120
transform 1 0 36616 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1607721120
transform 1 0 35328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1342_
timestamp 1607721120
transform 1 0 34868 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _0718_
timestamp 1607721120
transform 1 0 35420 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0713_
timestamp 1607721120
transform 1 0 36800 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_27_404
timestamp 1607721120
transform 1 0 38272 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_395
timestamp 1607721120
transform 1 0 37444 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_398
timestamp 1607721120
transform 1 0 37720 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_394
timestamp 1607721120
transform 1 0 37352 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1607721120
transform 1 0 38180 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1607721120
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1345_
timestamp 1607721120
transform 1 0 38456 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1344_
timestamp 1607721120
transform 1 0 37812 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_27_433
timestamp 1607721120
transform 1 0 40940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_425
timestamp 1607721120
transform 1 0 40204 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1607721120
transform 1 0 40940 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_418
timestamp 1607721120
transform 1 0 39560 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0707_
timestamp 1607721120
transform 1 0 40296 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_27_447
timestamp 1607721120
transform 1 0 42228 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_435
timestamp 1607721120
transform 1 0 41124 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1607721120
transform 1 0 42044 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1607721120
transform 1 0 41032 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_459
timestamp 1607721120
transform 1 0 43332 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_478
timestamp 1607721120
transform 1 0 45080 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_457
timestamp 1607721120
transform 1 0 43148 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1607721120
transform 1 0 43884 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1607721120
transform 1 0 43240 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1347_
timestamp 1607721120
transform 1 0 43976 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1346_
timestamp 1607721120
transform 1 0 43332 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_27_497
timestamp 1607721120
transform 1 0 46828 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_493
timestamp 1607721120
transform 1 0 46460 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_485
timestamp 1607721120
transform 1 0 45724 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1607721120
transform 1 0 46736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1348_
timestamp 1607721120
transform 1 0 45816 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_27_519
timestamp 1607721120
transform 1 0 48852 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_509
timestamp 1607721120
transform 1 0 47932 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_524
timestamp 1607721120
transform 1 0 49312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_520
timestamp 1607721120
transform 1 0 48944 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_517
timestamp 1607721120
transform 1 0 48668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_505
timestamp 1607721120
transform 1 0 47564 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1607721120
transform 1 0 48852 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1350_
timestamp 1607721120
transform 1 0 49404 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__or2_4  _0686_
timestamp 1607721120
transform 1 0 48208 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_27_547
timestamp 1607721120
transform 1 0 51428 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_535
timestamp 1607721120
transform 1 0 50324 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_544
timestamp 1607721120
transform 1 0 51152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1607721120
transform 1 0 49588 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0679_
timestamp 1607721120
transform 1 0 49680 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_27_559
timestamp 1607721120
transform 1 0 52532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_555
timestamp 1607721120
transform 1 0 52164 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_568
timestamp 1607721120
transform 1 0 53360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_556
timestamp 1607721120
transform 1 0 52256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1607721120
transform 1 0 52440 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_590
timestamp 1607721120
transform 1 0 55384 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_583
timestamp 1607721120
transform 1 0 54740 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_571
timestamp 1607721120
transform 1 0 53636 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_581
timestamp 1607721120
transform 1 0 54556 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1607721120
transform 1 0 55292 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1607721120
transform 1 0 54464 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1354_
timestamp 1607721120
transform 1 0 55292 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_27_614
timestamp 1607721120
transform 1 0 57592 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_602
timestamp 1607721120
transform 1 0 56488 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_608
timestamp 1607721120
transform 1 0 57040 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_633
timestamp 1607721120
transform 1 0 59340 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_621
timestamp 1607721120
transform 1 0 58236 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_632
timestamp 1607721120
transform 1 0 59248 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_620
timestamp 1607721120
transform 1 0 58144 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1607721120
transform 1 0 58144 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_645
timestamp 1607721120
transform 1 0 60444 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_640
timestamp 1607721120
transform 1 0 59984 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1607721120
transform 1 0 60076 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_660
timestamp 1607721120
transform 1 0 61824 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_652
timestamp 1607721120
transform 1 0 61088 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_660
timestamp 1607721120
transform 1 0 61824 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_654
timestamp 1607721120
transform 1 0 61272 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1607721120
transform 1 0 60996 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1607721120
transform -1 0 62192 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1607721120
transform -1 0 62192 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_642
timestamp 1607721120
transform 1 0 60168 0 -1 16864
box -38 -48 1142 592
<< labels >>
rlabel metal3 s 0 1096 800 1216 6 cen
port 0 nsew default tristate
rlabel metal3 s 0 3272 800 3392 6 set_out[0]
port 1 nsew default tristate
rlabel metal3 s 0 5448 800 5568 6 set_out[1]
port 2 nsew default tristate
rlabel metal3 s 0 7624 800 7744 6 set_out[2]
port 3 nsew default tristate
rlabel metal3 s 0 9800 800 9920 6 set_out[3]
port 4 nsew default tristate
rlabel metal3 s 0 11976 800 12096 6 shift_out[0]
port 5 nsew default tristate
rlabel metal3 s 0 14152 800 14272 6 shift_out[1]
port 6 nsew default tristate
rlabel metal3 s 0 16328 800 16448 6 shift_out[2]
port 7 nsew default tristate
rlabel metal3 s 0 18504 800 18624 6 shift_out[3]
port 8 nsew default tristate
rlabel metal2 s 386 0 442 800 6 wb_clk_i
port 9 nsew default input
rlabel metal2 s 1214 0 1270 800 6 wb_rst_i
port 10 nsew default input
rlabel metal2 s 938 18835 994 19635 6 wbs_ack_o
port 11 nsew default tristate
rlabel metal2 s 35898 0 35954 800 6 wbs_addr_i[0]
port 12 nsew default input
rlabel metal2 s 44546 0 44602 800 6 wbs_addr_i[10]
port 13 nsew default input
rlabel metal2 s 45466 0 45522 800 6 wbs_addr_i[11]
port 14 nsew default input
rlabel metal2 s 46294 0 46350 800 6 wbs_addr_i[12]
port 15 nsew default input
rlabel metal2 s 47122 0 47178 800 6 wbs_addr_i[13]
port 16 nsew default input
rlabel metal2 s 48042 0 48098 800 6 wbs_addr_i[14]
port 17 nsew default input
rlabel metal2 s 48870 0 48926 800 6 wbs_addr_i[15]
port 18 nsew default input
rlabel metal2 s 49790 0 49846 800 6 wbs_addr_i[16]
port 19 nsew default input
rlabel metal2 s 50618 0 50674 800 6 wbs_addr_i[17]
port 20 nsew default input
rlabel metal2 s 51538 0 51594 800 6 wbs_addr_i[18]
port 21 nsew default input
rlabel metal2 s 52366 0 52422 800 6 wbs_addr_i[19]
port 22 nsew default input
rlabel metal2 s 36726 0 36782 800 6 wbs_addr_i[1]
port 23 nsew default input
rlabel metal2 s 53194 0 53250 800 6 wbs_addr_i[20]
port 24 nsew default input
rlabel metal2 s 54114 0 54170 800 6 wbs_addr_i[21]
port 25 nsew default input
rlabel metal2 s 54942 0 54998 800 6 wbs_addr_i[22]
port 26 nsew default input
rlabel metal2 s 55862 0 55918 800 6 wbs_addr_i[23]
port 27 nsew default input
rlabel metal2 s 56690 0 56746 800 6 wbs_addr_i[24]
port 28 nsew default input
rlabel metal2 s 57610 0 57666 800 6 wbs_addr_i[25]
port 29 nsew default input
rlabel metal2 s 58438 0 58494 800 6 wbs_addr_i[26]
port 30 nsew default input
rlabel metal2 s 59266 0 59322 800 6 wbs_addr_i[27]
port 31 nsew default input
rlabel metal2 s 60186 0 60242 800 6 wbs_addr_i[28]
port 32 nsew default input
rlabel metal2 s 61014 0 61070 800 6 wbs_addr_i[29]
port 33 nsew default input
rlabel metal2 s 37646 0 37702 800 6 wbs_addr_i[2]
port 34 nsew default input
rlabel metal2 s 61934 0 61990 800 6 wbs_addr_i[30]
port 35 nsew default input
rlabel metal2 s 62762 0 62818 800 6 wbs_addr_i[31]
port 36 nsew default input
rlabel metal2 s 38474 0 38530 800 6 wbs_addr_i[3]
port 37 nsew default input
rlabel metal2 s 39394 0 39450 800 6 wbs_addr_i[4]
port 38 nsew default input
rlabel metal2 s 40222 0 40278 800 6 wbs_addr_i[5]
port 39 nsew default input
rlabel metal2 s 41050 0 41106 800 6 wbs_addr_i[6]
port 40 nsew default input
rlabel metal2 s 41970 0 42026 800 6 wbs_addr_i[7]
port 41 nsew default input
rlabel metal2 s 42798 0 42854 800 6 wbs_addr_i[8]
port 42 nsew default input
rlabel metal2 s 43718 0 43774 800 6 wbs_addr_i[9]
port 43 nsew default input
rlabel metal2 s 2962 0 3018 800 6 wbs_cyc_i
port 44 nsew default input
rlabel metal2 s 8114 0 8170 800 6 wbs_data_i[0]
port 45 nsew default input
rlabel metal2 s 16854 0 16910 800 6 wbs_data_i[10]
port 46 nsew default input
rlabel metal2 s 17682 0 17738 800 6 wbs_data_i[11]
port 47 nsew default input
rlabel metal2 s 18510 0 18566 800 6 wbs_data_i[12]
port 48 nsew default input
rlabel metal2 s 19430 0 19486 800 6 wbs_data_i[13]
port 49 nsew default input
rlabel metal2 s 20258 0 20314 800 6 wbs_data_i[14]
port 50 nsew default input
rlabel metal2 s 21178 0 21234 800 6 wbs_data_i[15]
port 51 nsew default input
rlabel metal2 s 22006 0 22062 800 6 wbs_data_i[16]
port 52 nsew default input
rlabel metal2 s 22926 0 22982 800 6 wbs_data_i[17]
port 53 nsew default input
rlabel metal2 s 23754 0 23810 800 6 wbs_data_i[18]
port 54 nsew default input
rlabel metal2 s 24582 0 24638 800 6 wbs_data_i[19]
port 55 nsew default input
rlabel metal2 s 9034 0 9090 800 6 wbs_data_i[1]
port 56 nsew default input
rlabel metal2 s 25502 0 25558 800 6 wbs_data_i[20]
port 57 nsew default input
rlabel metal2 s 26330 0 26386 800 6 wbs_data_i[21]
port 58 nsew default input
rlabel metal2 s 27250 0 27306 800 6 wbs_data_i[22]
port 59 nsew default input
rlabel metal2 s 28078 0 28134 800 6 wbs_data_i[23]
port 60 nsew default input
rlabel metal2 s 28998 0 29054 800 6 wbs_data_i[24]
port 61 nsew default input
rlabel metal2 s 29826 0 29882 800 6 wbs_data_i[25]
port 62 nsew default input
rlabel metal2 s 30654 0 30710 800 6 wbs_data_i[26]
port 63 nsew default input
rlabel metal2 s 31574 0 31630 800 6 wbs_data_i[27]
port 64 nsew default input
rlabel metal2 s 32402 0 32458 800 6 wbs_data_i[28]
port 65 nsew default input
rlabel metal2 s 33322 0 33378 800 6 wbs_data_i[29]
port 66 nsew default input
rlabel metal2 s 9862 0 9918 800 6 wbs_data_i[2]
port 67 nsew default input
rlabel metal2 s 34150 0 34206 800 6 wbs_data_i[30]
port 68 nsew default input
rlabel metal2 s 34978 0 35034 800 6 wbs_data_i[31]
port 69 nsew default input
rlabel metal2 s 10782 0 10838 800 6 wbs_data_i[3]
port 70 nsew default input
rlabel metal2 s 11610 0 11666 800 6 wbs_data_i[4]
port 71 nsew default input
rlabel metal2 s 12438 0 12494 800 6 wbs_data_i[5]
port 72 nsew default input
rlabel metal2 s 13358 0 13414 800 6 wbs_data_i[6]
port 73 nsew default input
rlabel metal2 s 14186 0 14242 800 6 wbs_data_i[7]
port 74 nsew default input
rlabel metal2 s 15106 0 15162 800 6 wbs_data_i[8]
port 75 nsew default input
rlabel metal2 s 15934 0 15990 800 6 wbs_data_i[9]
port 76 nsew default input
rlabel metal2 s 2778 18835 2834 19635 6 wbs_data_o[0]
port 77 nsew default tristate
rlabel metal2 s 22006 18835 22062 19635 6 wbs_data_o[10]
port 78 nsew default tristate
rlabel metal2 s 23938 18835 23994 19635 6 wbs_data_o[11]
port 79 nsew default tristate
rlabel metal2 s 25870 18835 25926 19635 6 wbs_data_o[12]
port 80 nsew default tristate
rlabel metal2 s 27710 18835 27766 19635 6 wbs_data_o[13]
port 81 nsew default tristate
rlabel metal2 s 29642 18835 29698 19635 6 wbs_data_o[14]
port 82 nsew default tristate
rlabel metal2 s 31574 18835 31630 19635 6 wbs_data_o[15]
port 83 nsew default tristate
rlabel metal2 s 33506 18835 33562 19635 6 wbs_data_o[16]
port 84 nsew default tristate
rlabel metal2 s 35438 18835 35494 19635 6 wbs_data_o[17]
port 85 nsew default tristate
rlabel metal2 s 37370 18835 37426 19635 6 wbs_data_o[18]
port 86 nsew default tristate
rlabel metal2 s 39210 18835 39266 19635 6 wbs_data_o[19]
port 87 nsew default tristate
rlabel metal2 s 4710 18835 4766 19635 6 wbs_data_o[1]
port 88 nsew default tristate
rlabel metal2 s 41142 18835 41198 19635 6 wbs_data_o[20]
port 89 nsew default tristate
rlabel metal2 s 43074 18835 43130 19635 6 wbs_data_o[21]
port 90 nsew default tristate
rlabel metal2 s 45006 18835 45062 19635 6 wbs_data_o[22]
port 91 nsew default tristate
rlabel metal2 s 46938 18835 46994 19635 6 wbs_data_o[23]
port 92 nsew default tristate
rlabel metal2 s 48870 18835 48926 19635 6 wbs_data_o[24]
port 93 nsew default tristate
rlabel metal2 s 50802 18835 50858 19635 6 wbs_data_o[25]
port 94 nsew default tristate
rlabel metal2 s 52642 18835 52698 19635 6 wbs_data_o[26]
port 95 nsew default tristate
rlabel metal2 s 54574 18835 54630 19635 6 wbs_data_o[27]
port 96 nsew default tristate
rlabel metal2 s 56506 18835 56562 19635 6 wbs_data_o[28]
port 97 nsew default tristate
rlabel metal2 s 58438 18835 58494 19635 6 wbs_data_o[29]
port 98 nsew default tristate
rlabel metal2 s 6642 18835 6698 19635 6 wbs_data_o[2]
port 99 nsew default tristate
rlabel metal2 s 60370 18835 60426 19635 6 wbs_data_o[30]
port 100 nsew default tristate
rlabel metal2 s 62302 18835 62358 19635 6 wbs_data_o[31]
port 101 nsew default tristate
rlabel metal2 s 8574 18835 8630 19635 6 wbs_data_o[3]
port 102 nsew default tristate
rlabel metal2 s 10506 18835 10562 19635 6 wbs_data_o[4]
port 103 nsew default tristate
rlabel metal2 s 12438 18835 12494 19635 6 wbs_data_o[5]
port 104 nsew default tristate
rlabel metal2 s 14278 18835 14334 19635 6 wbs_data_o[6]
port 105 nsew default tristate
rlabel metal2 s 16210 18835 16266 19635 6 wbs_data_o[7]
port 106 nsew default tristate
rlabel metal2 s 18142 18835 18198 19635 6 wbs_data_o[8]
port 107 nsew default tristate
rlabel metal2 s 20074 18835 20130 19635 6 wbs_data_o[9]
port 108 nsew default tristate
rlabel metal2 s 4710 0 4766 800 6 wbs_sel_i[0]
port 109 nsew default input
rlabel metal2 s 5538 0 5594 800 6 wbs_sel_i[1]
port 110 nsew default input
rlabel metal2 s 6366 0 6422 800 6 wbs_sel_i[2]
port 111 nsew default input
rlabel metal2 s 7286 0 7342 800 6 wbs_sel_i[3]
port 112 nsew default input
rlabel metal2 s 2042 0 2098 800 6 wbs_stb_i
port 113 nsew default input
rlabel metal2 s 3790 0 3846 800 6 wbs_we_i
port 114 nsew default input
rlabel metal4 s 11125 2128 11445 17456 6 VPWR
port 115 nsew default input
rlabel metal4 s 21307 2128 21627 17456 6 VGND
port 116 nsew default input
<< properties >>
string FIXED_BBOX 0 0 62822 19635
<< end >>

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 3198.900 BY 3888.080 ;
  PIN gpio_east[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 75.440 3149.480 76.040 ;
    END
  END gpio_east[0]
  PIN gpio_east[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 138.680 3149.480 139.280 ;
    END
  END gpio_east[1]
  PIN gpio_east[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 201.920 3149.480 202.520 ;
    END
  END gpio_east[2]
  PIN gpio_east[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 265.160 3149.480 265.760 ;
    END
  END gpio_east[3]
  PIN gpio_east[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 328.400 3149.480 329.000 ;
    END
  END gpio_east[4]
  PIN gpio_east[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 391.640 3149.480 392.240 ;
    END
  END gpio_east[5]
  PIN gpio_east[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 454.880 3149.480 455.480 ;
    END
  END gpio_east[6]
  PIN gpio_east[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 518.120 3149.480 518.720 ;
    END
  END gpio_east[7]
  PIN gpio_east[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 582.040 3149.480 582.640 ;
    END
  END gpio_east[8]
  PIN gpio_east[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 645.280 3149.480 645.880 ;
    END
  END gpio_east[9]
  PIN gpio_north[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 93.730 3840.120 94.010 3844.120 ;
    END
  END gpio_north[0]
  PIN gpio_north[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 182.050 3840.120 182.330 3844.120 ;
    END
  END gpio_north[1]
  PIN gpio_north[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 270.830 3840.120 271.110 3844.120 ;
    END
  END gpio_north[2]
  PIN gpio_north[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 359.150 3840.120 359.430 3844.120 ;
    END
  END gpio_north[3]
  PIN gpio_north[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 447.930 3840.120 448.210 3844.120 ;
    END
  END gpio_north[4]
  PIN gpio_north[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 536.250 3840.120 536.530 3844.120 ;
    END
  END gpio_north[5]
  PIN gpio_north[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 625.030 3840.120 625.310 3844.120 ;
    END
  END gpio_north[6]
  PIN gpio_north[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 713.350 3840.120 713.630 3844.120 ;
    END
  END gpio_north[7]
  PIN gpio_north[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 802.130 3840.120 802.410 3844.120 ;
    END
  END gpio_north[8]
  PIN gpio_north[9]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 890.450 3840.120 890.730 3844.120 ;
    END
  END gpio_north[9]
  PIN gpio_south[0]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 111.210 44.120 111.490 48.120 ;
    END
  END gpio_south[0]
  PIN gpio_south[1]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 234.950 44.120 235.230 48.120 ;
    END
  END gpio_south[1]
  PIN gpio_south[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 359.150 44.120 359.430 48.120 ;
    END
  END gpio_south[2]
  PIN gpio_south[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 482.890 44.120 483.170 48.120 ;
    END
  END gpio_south[3]
  PIN gpio_south[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 607.090 44.120 607.370 48.120 ;
    END
  END gpio_south[4]
  PIN gpio_south[5]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 730.830 44.120 731.110 48.120 ;
    END
  END gpio_south[5]
  PIN gpio_south[6]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 855.030 44.120 855.310 48.120 ;
    END
  END gpio_south[6]
  PIN gpio_south[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 978.770 44.120 979.050 48.120 ;
    END
  END gpio_south[7]
  PIN gpio_west[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 123.040 53.480 123.640 ;
    END
  END gpio_west[0]
  PIN gpio_west[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 280.800 53.480 281.400 ;
    END
  END gpio_west[1]
  PIN gpio_west[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 439.240 53.480 439.840 ;
    END
  END gpio_west[2]
  PIN gpio_west[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 597.680 53.480 598.280 ;
    END
  END gpio_west[3]
  PIN gpio_west[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 756.120 53.480 756.720 ;
    END
  END gpio_west[4]
  PIN gpio_west[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 914.560 53.480 915.160 ;
    END
  END gpio_west[5]
  PIN gpio_west[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1073.000 53.480 1073.600 ;
    END
  END gpio_west[6]
  PIN gpio_west[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1230.760 53.480 1231.360 ;
    END
  END gpio_west[7]
  PIN gpio_west[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1389.200 53.480 1389.800 ;
    END
  END gpio_west[8]
  PIN gpio_west[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1547.640 53.480 1548.240 ;
    END
  END gpio_west[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2734.920 3149.480 2735.520 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2798.160 3149.480 2798.760 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.970 44.120 1103.250 48.120 ;
    END
  END wbs_ack_o
  PIN wbs_addr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 979.230 3840.120 979.510 3844.120 ;
    END
  END wbs_addr_i[0]
  PIN wbs_addr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1245.110 3840.120 1245.390 3844.120 ;
    END
  END wbs_addr_i[10]
  PIN wbs_addr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1598.850 44.120 1599.130 48.120 ;
    END
  END wbs_addr_i[11]
  PIN wbs_addr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1333.430 3840.120 1333.710 3844.120 ;
    END
  END wbs_addr_i[12]
  PIN wbs_addr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1422.210 3840.120 1422.490 3844.120 ;
    END
  END wbs_addr_i[13]
  PIN wbs_addr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1510.530 3840.120 1510.810 3844.120 ;
    END
  END wbs_addr_i[14]
  PIN wbs_addr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1864.520 53.480 1865.120 ;
    END
  END wbs_addr_i[15]
  PIN wbs_addr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 3051.800 3149.480 3052.400 ;
    END
  END wbs_addr_i[16]
  PIN wbs_addr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2022.960 53.480 2023.560 ;
    END
  END wbs_addr_i[17]
  PIN wbs_addr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 3115.040 3149.480 3115.640 ;
    END
  END wbs_addr_i[18]
  PIN wbs_addr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2180.720 53.480 2181.320 ;
    END
  END wbs_addr_i[19]
  PIN wbs_addr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 1706.080 53.480 1706.680 ;
    END
  END wbs_addr_i[1]
  PIN wbs_addr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1599.310 3840.120 1599.590 3844.120 ;
    END
  END wbs_addr_i[20]
  PIN wbs_addr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1687.630 3840.120 1687.910 3844.120 ;
    END
  END wbs_addr_i[21]
  PIN wbs_addr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1776.410 3840.120 1776.690 3844.120 ;
    END
  END wbs_addr_i[22]
  PIN wbs_addr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1723.050 44.120 1723.330 48.120 ;
    END
  END wbs_addr_i[23]
  PIN wbs_addr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1864.730 3840.120 1865.010 3844.120 ;
    END
  END wbs_addr_i[24]
  PIN wbs_addr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1846.790 44.120 1847.070 48.120 ;
    END
  END wbs_addr_i[25]
  PIN wbs_addr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.510 3840.120 1953.790 3844.120 ;
    END
  END wbs_addr_i[26]
  PIN wbs_addr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 3178.280 3149.480 3178.880 ;
    END
  END wbs_addr_i[27]
  PIN wbs_addr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2339.160 53.480 2339.760 ;
    END
  END wbs_addr_i[28]
  PIN wbs_addr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2497.600 53.480 2498.200 ;
    END
  END wbs_addr_i[29]
  PIN wbs_addr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2861.400 3149.480 2862.000 ;
    END
  END wbs_addr_i[2]
  PIN wbs_addr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1970.990 44.120 1971.270 48.120 ;
    END
  END wbs_addr_i[30]
  PIN wbs_addr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 3241.520 3149.480 3242.120 ;
    END
  END wbs_addr_i[31]
  PIN wbs_addr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1067.550 3840.120 1067.830 3844.120 ;
    END
  END wbs_addr_i[3]
  PIN wbs_addr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1227.170 44.120 1227.450 48.120 ;
    END
  END wbs_addr_i[4]
  PIN wbs_addr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1350.910 44.120 1351.190 48.120 ;
    END
  END wbs_addr_i[5]
  PIN wbs_addr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2925.320 3149.480 2925.920 ;
    END
  END wbs_addr_i[6]
  PIN wbs_addr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1156.330 3840.120 1156.610 3844.120 ;
    END
  END wbs_addr_i[7]
  PIN wbs_addr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2988.560 3149.480 2989.160 ;
    END
  END wbs_addr_i[8]
  PIN wbs_addr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1475.110 44.120 1475.390 48.120 ;
    END
  END wbs_addr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2094.730 44.120 2095.010 48.120 ;
    END
  END wbs_cyc_i
  PIN wbs_data_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2041.830 3840.120 2042.110 3844.120 ;
    END
  END wbs_data_i[0]
  PIN wbs_data_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2396.490 3840.120 2396.770 3844.120 ;
    END
  END wbs_data_i[10]
  PIN wbs_data_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2814.480 53.480 2815.080 ;
    END
  END wbs_data_i[11]
  PIN wbs_data_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 3431.920 3149.480 3432.520 ;
    END
  END wbs_data_i[12]
  PIN wbs_data_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2972.920 53.480 2973.520 ;
    END
  END wbs_data_i[13]
  PIN wbs_data_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 3495.160 3149.480 3495.760 ;
    END
  END wbs_data_i[14]
  PIN wbs_data_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 3558.400 3149.480 3559.000 ;
    END
  END wbs_data_i[15]
  PIN wbs_data_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2484.810 3840.120 2485.090 3844.120 ;
    END
  END wbs_data_i[16]
  PIN wbs_data_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2573.590 3840.120 2573.870 3844.120 ;
    END
  END wbs_data_i[17]
  PIN wbs_data_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.910 3840.120 2662.190 3844.120 ;
    END
  END wbs_data_i[18]
  PIN wbs_data_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3130.680 53.480 3131.280 ;
    END
  END wbs_data_i[19]
  PIN wbs_data_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 2656.040 53.480 2656.640 ;
    END
  END wbs_data_i[1]
  PIN wbs_data_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 3621.640 3149.480 3622.240 ;
    END
  END wbs_data_i[20]
  PIN wbs_data_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2591.070 44.120 2591.350 48.120 ;
    END
  END wbs_data_i[21]
  PIN wbs_data_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3289.120 53.480 3289.720 ;
    END
  END wbs_data_i[22]
  PIN wbs_data_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3447.560 53.480 3448.160 ;
    END
  END wbs_data_i[23]
  PIN wbs_data_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.810 44.120 2715.090 48.120 ;
    END
  END wbs_data_i[24]
  PIN wbs_data_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3606.000 53.480 3606.600 ;
    END
  END wbs_data_i[25]
  PIN wbs_data_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.010 44.120 2839.290 48.120 ;
    END
  END wbs_data_i[26]
  PIN wbs_data_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.690 3840.120 2750.970 3844.120 ;
    END
  END wbs_data_i[27]
  PIN wbs_data_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2962.750 44.120 2963.030 48.120 ;
    END
  END wbs_data_i[28]
  PIN wbs_data_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.010 3840.120 2839.290 3844.120 ;
    END
  END wbs_data_i[29]
  PIN wbs_data_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2130.610 3840.120 2130.890 3844.120 ;
    END
  END wbs_data_i[2]
  PIN wbs_data_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3086.950 44.120 3087.230 48.120 ;
    END
  END wbs_data_i[30]
  PIN wbs_data_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2927.790 3840.120 2928.070 3844.120 ;
    END
  END wbs_data_i[31]
  PIN wbs_data_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 3304.760 3149.480 3305.360 ;
    END
  END wbs_data_i[3]
  PIN wbs_data_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2218.930 44.120 2219.210 48.120 ;
    END
  END wbs_data_i[4]
  PIN wbs_data_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2343.130 44.120 2343.410 48.120 ;
    END
  END wbs_data_i[5]
  PIN wbs_data_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2219.390 3840.120 2219.670 3844.120 ;
    END
  END wbs_data_i[6]
  PIN wbs_data_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2307.710 3840.120 2307.990 3844.120 ;
    END
  END wbs_data_i[7]
  PIN wbs_data_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2466.870 44.120 2467.150 48.120 ;
    END
  END wbs_data_i[8]
  PIN wbs_data_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 3368.000 3149.480 3368.600 ;
    END
  END wbs_data_i[9]
  PIN wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 708.520 3149.480 709.120 ;
    END
  END wbs_data_o[0]
  PIN wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1341.600 3149.480 1342.200 ;
    END
  END wbs_data_o[10]
  PIN wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1404.840 3149.480 1405.440 ;
    END
  END wbs_data_o[11]
  PIN wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1468.080 3149.480 1468.680 ;
    END
  END wbs_data_o[12]
  PIN wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1532.000 3149.480 1532.600 ;
    END
  END wbs_data_o[13]
  PIN wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1595.240 3149.480 1595.840 ;
    END
  END wbs_data_o[14]
  PIN wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1658.480 3149.480 1659.080 ;
    END
  END wbs_data_o[15]
  PIN wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1721.720 3149.480 1722.320 ;
    END
  END wbs_data_o[16]
  PIN wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1784.960 3149.480 1785.560 ;
    END
  END wbs_data_o[17]
  PIN wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1848.200 3149.480 1848.800 ;
    END
  END wbs_data_o[18]
  PIN wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1911.440 3149.480 1912.040 ;
    END
  END wbs_data_o[19]
  PIN wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 771.760 3149.480 772.360 ;
    END
  END wbs_data_o[1]
  PIN wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1975.360 3149.480 1975.960 ;
    END
  END wbs_data_o[20]
  PIN wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2038.600 3149.480 2039.200 ;
    END
  END wbs_data_o[21]
  PIN wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2101.840 3149.480 2102.440 ;
    END
  END wbs_data_o[22]
  PIN wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2165.080 3149.480 2165.680 ;
    END
  END wbs_data_o[23]
  PIN wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2228.320 3149.480 2228.920 ;
    END
  END wbs_data_o[24]
  PIN wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2291.560 3149.480 2292.160 ;
    END
  END wbs_data_o[25]
  PIN wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2354.800 3149.480 2355.400 ;
    END
  END wbs_data_o[26]
  PIN wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2418.040 3149.480 2418.640 ;
    END
  END wbs_data_o[27]
  PIN wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2481.960 3149.480 2482.560 ;
    END
  END wbs_data_o[28]
  PIN wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2545.200 3149.480 2545.800 ;
    END
  END wbs_data_o[29]
  PIN wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 835.000 3149.480 835.600 ;
    END
  END wbs_data_o[2]
  PIN wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2608.440 3149.480 2609.040 ;
    END
  END wbs_data_o[30]
  PIN wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 2671.680 3149.480 2672.280 ;
    END
  END wbs_data_o[31]
  PIN wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 898.240 3149.480 898.840 ;
    END
  END wbs_data_o[3]
  PIN wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 961.480 3149.480 962.080 ;
    END
  END wbs_data_o[4]
  PIN wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1025.400 3149.480 1026.000 ;
    END
  END wbs_data_o[5]
  PIN wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1088.640 3149.480 1089.240 ;
    END
  END wbs_data_o[6]
  PIN wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1151.880 3149.480 1152.480 ;
    END
  END wbs_data_o[7]
  PIN wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1215.120 3149.480 1215.720 ;
    END
  END wbs_data_o[8]
  PIN wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 3145.480 1278.360 3149.480 1278.960 ;
    END
  END wbs_data_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3016.110 3840.120 3016.390 3844.120 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 3684.880 3149.480 3685.480 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3104.890 3840.120 3105.170 3844.120 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 3764.440 53.480 3765.040 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 3748.120 3149.480 3748.720 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 3145.480 3811.360 3149.480 3811.960 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 25.000 25.000 3173.900 45.000 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.000 3198.900 20.000 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 55.000 54.915 3143.900 3833.165 ;
      LAYER met1 ;
        RECT 55.000 54.760 3143.900 3833.320 ;
      LAYER met2 ;
        RECT 63.370 3839.840 93.450 3840.120 ;
        RECT 94.290 3839.840 181.770 3840.120 ;
        RECT 182.610 3839.840 270.550 3840.120 ;
        RECT 271.390 3839.840 358.870 3840.120 ;
        RECT 359.710 3839.840 447.650 3840.120 ;
        RECT 448.490 3839.840 535.970 3840.120 ;
        RECT 536.810 3839.840 624.750 3840.120 ;
        RECT 625.590 3839.840 713.070 3840.120 ;
        RECT 713.910 3839.840 801.850 3840.120 ;
        RECT 802.690 3839.840 890.170 3840.120 ;
        RECT 891.010 3839.840 978.950 3840.120 ;
        RECT 979.790 3839.840 1067.270 3840.120 ;
        RECT 1068.110 3839.840 1156.050 3840.120 ;
        RECT 1156.890 3839.840 1244.830 3840.120 ;
        RECT 1245.670 3839.840 1333.150 3840.120 ;
        RECT 1333.990 3839.840 1421.930 3840.120 ;
        RECT 1422.770 3839.840 1510.250 3840.120 ;
        RECT 1511.090 3839.840 1599.030 3840.120 ;
        RECT 1599.870 3839.840 1687.350 3840.120 ;
        RECT 1688.190 3839.840 1776.130 3840.120 ;
        RECT 1776.970 3839.840 1864.450 3840.120 ;
        RECT 1865.290 3839.840 1953.230 3840.120 ;
        RECT 1954.070 3839.840 2041.550 3840.120 ;
        RECT 2042.390 3839.840 2130.330 3840.120 ;
        RECT 2131.170 3839.840 2219.110 3840.120 ;
        RECT 2219.950 3839.840 2307.430 3840.120 ;
        RECT 2308.270 3839.840 2396.210 3840.120 ;
        RECT 2397.050 3839.840 2484.530 3840.120 ;
        RECT 2485.370 3839.840 2573.310 3840.120 ;
        RECT 2574.150 3839.840 2661.630 3840.120 ;
        RECT 2662.470 3839.840 2750.410 3840.120 ;
        RECT 2751.250 3839.840 2838.730 3840.120 ;
        RECT 2839.570 3839.840 2927.510 3840.120 ;
        RECT 2928.350 3839.840 3015.830 3840.120 ;
        RECT 3016.670 3839.840 3104.610 3840.120 ;
        RECT 3105.450 3839.840 3133.690 3840.120 ;
        RECT 63.370 48.400 3133.690 3839.840 ;
        RECT 63.370 48.120 110.930 48.400 ;
        RECT 111.770 48.120 234.670 48.400 ;
        RECT 235.510 48.120 358.870 48.400 ;
        RECT 359.710 48.120 482.610 48.400 ;
        RECT 483.450 48.120 606.810 48.400 ;
        RECT 607.650 48.120 730.550 48.400 ;
        RECT 731.390 48.120 854.750 48.400 ;
        RECT 855.590 48.120 978.490 48.400 ;
        RECT 979.330 48.120 1102.690 48.400 ;
        RECT 1103.530 48.120 1226.890 48.400 ;
        RECT 1227.730 48.120 1350.630 48.400 ;
        RECT 1351.470 48.120 1474.830 48.400 ;
        RECT 1475.670 48.120 1598.570 48.400 ;
        RECT 1599.410 48.120 1722.770 48.400 ;
        RECT 1723.610 48.120 1846.510 48.400 ;
        RECT 1847.350 48.120 1970.710 48.400 ;
        RECT 1971.550 48.120 2094.450 48.400 ;
        RECT 2095.290 48.120 2218.650 48.400 ;
        RECT 2219.490 48.120 2342.850 48.400 ;
        RECT 2343.690 48.120 2466.590 48.400 ;
        RECT 2467.430 48.120 2590.790 48.400 ;
        RECT 2591.630 48.120 2714.530 48.400 ;
        RECT 2715.370 48.120 2838.730 48.400 ;
        RECT 2839.570 48.120 2962.470 48.400 ;
        RECT 2963.310 48.120 3086.670 48.400 ;
        RECT 3087.510 48.120 3133.690 48.400 ;
      LAYER met3 ;
        RECT 53.480 3812.360 3145.480 3833.245 ;
        RECT 53.480 3810.960 3145.080 3812.360 ;
        RECT 53.480 3765.440 3145.480 3810.960 ;
        RECT 53.880 3764.040 3145.480 3765.440 ;
        RECT 53.480 3749.120 3145.480 3764.040 ;
        RECT 53.480 3747.720 3145.080 3749.120 ;
        RECT 53.480 3685.880 3145.480 3747.720 ;
        RECT 53.480 3684.480 3145.080 3685.880 ;
        RECT 53.480 3622.640 3145.480 3684.480 ;
        RECT 53.480 3621.240 3145.080 3622.640 ;
        RECT 53.480 3607.000 3145.480 3621.240 ;
        RECT 53.880 3605.600 3145.480 3607.000 ;
        RECT 53.480 3559.400 3145.480 3605.600 ;
        RECT 53.480 3558.000 3145.080 3559.400 ;
        RECT 53.480 3496.160 3145.480 3558.000 ;
        RECT 53.480 3494.760 3145.080 3496.160 ;
        RECT 53.480 3448.560 3145.480 3494.760 ;
        RECT 53.880 3447.160 3145.480 3448.560 ;
        RECT 53.480 3432.920 3145.480 3447.160 ;
        RECT 53.480 3431.520 3145.080 3432.920 ;
        RECT 53.480 3369.000 3145.480 3431.520 ;
        RECT 53.480 3367.600 3145.080 3369.000 ;
        RECT 53.480 3305.760 3145.480 3367.600 ;
        RECT 53.480 3304.360 3145.080 3305.760 ;
        RECT 53.480 3290.120 3145.480 3304.360 ;
        RECT 53.880 3288.720 3145.480 3290.120 ;
        RECT 53.480 3242.520 3145.480 3288.720 ;
        RECT 53.480 3241.120 3145.080 3242.520 ;
        RECT 53.480 3179.280 3145.480 3241.120 ;
        RECT 53.480 3177.880 3145.080 3179.280 ;
        RECT 53.480 3131.680 3145.480 3177.880 ;
        RECT 53.880 3130.280 3145.480 3131.680 ;
        RECT 53.480 3116.040 3145.480 3130.280 ;
        RECT 53.480 3114.640 3145.080 3116.040 ;
        RECT 53.480 3052.800 3145.480 3114.640 ;
        RECT 53.480 3051.400 3145.080 3052.800 ;
        RECT 53.480 2989.560 3145.480 3051.400 ;
        RECT 53.480 2988.160 3145.080 2989.560 ;
        RECT 53.480 2973.920 3145.480 2988.160 ;
        RECT 53.880 2972.520 3145.480 2973.920 ;
        RECT 53.480 2926.320 3145.480 2972.520 ;
        RECT 53.480 2924.920 3145.080 2926.320 ;
        RECT 53.480 2862.400 3145.480 2924.920 ;
        RECT 53.480 2861.000 3145.080 2862.400 ;
        RECT 53.480 2815.480 3145.480 2861.000 ;
        RECT 53.880 2814.080 3145.480 2815.480 ;
        RECT 53.480 2799.160 3145.480 2814.080 ;
        RECT 53.480 2797.760 3145.080 2799.160 ;
        RECT 53.480 2735.920 3145.480 2797.760 ;
        RECT 53.480 2734.520 3145.080 2735.920 ;
        RECT 53.480 2672.680 3145.480 2734.520 ;
        RECT 53.480 2671.280 3145.080 2672.680 ;
        RECT 53.480 2657.040 3145.480 2671.280 ;
        RECT 53.880 2655.640 3145.480 2657.040 ;
        RECT 53.480 2609.440 3145.480 2655.640 ;
        RECT 53.480 2608.040 3145.080 2609.440 ;
        RECT 53.480 2546.200 3145.480 2608.040 ;
        RECT 53.480 2544.800 3145.080 2546.200 ;
        RECT 53.480 2498.600 3145.480 2544.800 ;
        RECT 53.880 2497.200 3145.480 2498.600 ;
        RECT 53.480 2482.960 3145.480 2497.200 ;
        RECT 53.480 2481.560 3145.080 2482.960 ;
        RECT 53.480 2419.040 3145.480 2481.560 ;
        RECT 53.480 2417.640 3145.080 2419.040 ;
        RECT 53.480 2355.800 3145.480 2417.640 ;
        RECT 53.480 2354.400 3145.080 2355.800 ;
        RECT 53.480 2340.160 3145.480 2354.400 ;
        RECT 53.880 2338.760 3145.480 2340.160 ;
        RECT 53.480 2292.560 3145.480 2338.760 ;
        RECT 53.480 2291.160 3145.080 2292.560 ;
        RECT 53.480 2229.320 3145.480 2291.160 ;
        RECT 53.480 2227.920 3145.080 2229.320 ;
        RECT 53.480 2181.720 3145.480 2227.920 ;
        RECT 53.880 2180.320 3145.480 2181.720 ;
        RECT 53.480 2166.080 3145.480 2180.320 ;
        RECT 53.480 2164.680 3145.080 2166.080 ;
        RECT 53.480 2102.840 3145.480 2164.680 ;
        RECT 53.480 2101.440 3145.080 2102.840 ;
        RECT 53.480 2039.600 3145.480 2101.440 ;
        RECT 53.480 2038.200 3145.080 2039.600 ;
        RECT 53.480 2023.960 3145.480 2038.200 ;
        RECT 53.880 2022.560 3145.480 2023.960 ;
        RECT 53.480 1976.360 3145.480 2022.560 ;
        RECT 53.480 1974.960 3145.080 1976.360 ;
        RECT 53.480 1912.440 3145.480 1974.960 ;
        RECT 53.480 1911.040 3145.080 1912.440 ;
        RECT 53.480 1865.520 3145.480 1911.040 ;
        RECT 53.880 1864.120 3145.480 1865.520 ;
        RECT 53.480 1849.200 3145.480 1864.120 ;
        RECT 53.480 1847.800 3145.080 1849.200 ;
        RECT 53.480 1785.960 3145.480 1847.800 ;
        RECT 53.480 1784.560 3145.080 1785.960 ;
        RECT 53.480 1722.720 3145.480 1784.560 ;
        RECT 53.480 1721.320 3145.080 1722.720 ;
        RECT 53.480 1707.080 3145.480 1721.320 ;
        RECT 53.880 1705.680 3145.480 1707.080 ;
        RECT 53.480 1659.480 3145.480 1705.680 ;
        RECT 53.480 1658.080 3145.080 1659.480 ;
        RECT 53.480 1596.240 3145.480 1658.080 ;
        RECT 53.480 1594.840 3145.080 1596.240 ;
        RECT 53.480 1548.640 3145.480 1594.840 ;
        RECT 53.880 1547.240 3145.480 1548.640 ;
        RECT 53.480 1533.000 3145.480 1547.240 ;
        RECT 53.480 1531.600 3145.080 1533.000 ;
        RECT 53.480 1469.080 3145.480 1531.600 ;
        RECT 53.480 1467.680 3145.080 1469.080 ;
        RECT 53.480 1405.840 3145.480 1467.680 ;
        RECT 53.480 1404.440 3145.080 1405.840 ;
        RECT 53.480 1390.200 3145.480 1404.440 ;
        RECT 53.880 1388.800 3145.480 1390.200 ;
        RECT 53.480 1342.600 3145.480 1388.800 ;
        RECT 53.480 1341.200 3145.080 1342.600 ;
        RECT 53.480 1279.360 3145.480 1341.200 ;
        RECT 53.480 1277.960 3145.080 1279.360 ;
        RECT 53.480 1231.760 3145.480 1277.960 ;
        RECT 53.880 1230.360 3145.480 1231.760 ;
        RECT 53.480 1216.120 3145.480 1230.360 ;
        RECT 53.480 1214.720 3145.080 1216.120 ;
        RECT 53.480 1152.880 3145.480 1214.720 ;
        RECT 53.480 1151.480 3145.080 1152.880 ;
        RECT 53.480 1089.640 3145.480 1151.480 ;
        RECT 53.480 1088.240 3145.080 1089.640 ;
        RECT 53.480 1074.000 3145.480 1088.240 ;
        RECT 53.880 1072.600 3145.480 1074.000 ;
        RECT 53.480 1026.400 3145.480 1072.600 ;
        RECT 53.480 1025.000 3145.080 1026.400 ;
        RECT 53.480 962.480 3145.480 1025.000 ;
        RECT 53.480 961.080 3145.080 962.480 ;
        RECT 53.480 915.560 3145.480 961.080 ;
        RECT 53.880 914.160 3145.480 915.560 ;
        RECT 53.480 899.240 3145.480 914.160 ;
        RECT 53.480 897.840 3145.080 899.240 ;
        RECT 53.480 836.000 3145.480 897.840 ;
        RECT 53.480 834.600 3145.080 836.000 ;
        RECT 53.480 772.760 3145.480 834.600 ;
        RECT 53.480 771.360 3145.080 772.760 ;
        RECT 53.480 757.120 3145.480 771.360 ;
        RECT 53.880 755.720 3145.480 757.120 ;
        RECT 53.480 709.520 3145.480 755.720 ;
        RECT 53.480 708.120 3145.080 709.520 ;
        RECT 53.480 646.280 3145.480 708.120 ;
        RECT 53.480 644.880 3145.080 646.280 ;
        RECT 53.480 598.680 3145.480 644.880 ;
        RECT 53.880 597.280 3145.480 598.680 ;
        RECT 53.480 583.040 3145.480 597.280 ;
        RECT 53.480 581.640 3145.080 583.040 ;
        RECT 53.480 519.120 3145.480 581.640 ;
        RECT 53.480 517.720 3145.080 519.120 ;
        RECT 53.480 455.880 3145.480 517.720 ;
        RECT 53.480 454.480 3145.080 455.880 ;
        RECT 53.480 440.240 3145.480 454.480 ;
        RECT 53.880 438.840 3145.480 440.240 ;
        RECT 53.480 392.640 3145.480 438.840 ;
        RECT 53.480 391.240 3145.080 392.640 ;
        RECT 53.480 329.400 3145.480 391.240 ;
        RECT 53.480 328.000 3145.080 329.400 ;
        RECT 53.480 281.800 3145.480 328.000 ;
        RECT 53.880 280.400 3145.480 281.800 ;
        RECT 53.480 266.160 3145.480 280.400 ;
        RECT 53.480 264.760 3145.080 266.160 ;
        RECT 53.480 202.920 3145.480 264.760 ;
        RECT 53.480 201.520 3145.080 202.920 ;
        RECT 53.480 139.680 3145.480 201.520 ;
        RECT 53.480 138.280 3145.080 139.680 ;
        RECT 53.480 124.040 3145.480 138.280 ;
        RECT 53.880 122.640 3145.480 124.040 ;
        RECT 53.480 76.440 3145.480 122.640 ;
        RECT 53.480 75.040 3145.080 76.440 ;
        RECT 53.480 54.835 3145.480 75.040 ;
      LAYER met4 ;
        RECT 0.000 0.000 3198.900 3888.080 ;
      LAYER met5 ;
        RECT 0.000 70.610 3198.900 3888.080 ;
  END
END fpga
END LIBRARY


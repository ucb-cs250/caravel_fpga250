VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.090 92.635 2898.370 93.005 ;
        RECT 2898.160 88.245 2898.300 92.635 ;
        RECT 2898.090 87.875 2898.370 88.245 ;
      LAYER via2 ;
        RECT 2898.090 92.680 2898.370 92.960 ;
        RECT 2898.090 87.920 2898.370 88.200 ;
      LAYER met3 ;
        RECT 2881.000 95.560 2885.000 96.160 ;
        RECT 2884.510 92.970 2884.810 95.560 ;
        RECT 2898.065 92.970 2898.395 92.985 ;
        RECT 2884.510 92.670 2898.395 92.970 ;
        RECT 2898.065 92.655 2898.395 92.670 ;
        RECT 2898.065 88.210 2898.395 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.065 87.910 2924.800 88.210 ;
        RECT 2898.065 87.895 2898.395 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1037.370 3445.460 1037.690 3445.520 ;
        RECT 2880.590 3445.460 2880.910 3445.520 ;
        RECT 1037.370 3445.320 2880.910 3445.460 ;
        RECT 1037.370 3445.260 1037.690 3445.320 ;
        RECT 2880.590 3445.260 2880.910 3445.320 ;
        RECT 2880.590 2435.660 2880.910 2435.720 ;
        RECT 2898.530 2435.660 2898.850 2435.720 ;
        RECT 2880.590 2435.520 2898.850 2435.660 ;
        RECT 2880.590 2435.460 2880.910 2435.520 ;
        RECT 2898.530 2435.460 2898.850 2435.520 ;
      LAYER via ;
        RECT 1037.400 3445.260 1037.660 3445.520 ;
        RECT 2880.620 3445.260 2880.880 3445.520 ;
        RECT 2880.620 2435.460 2880.880 2435.720 ;
        RECT 2898.560 2435.460 2898.820 2435.720 ;
      LAYER met2 ;
        RECT 1037.400 3445.230 1037.660 3445.550 ;
        RECT 2880.620 3445.230 2880.880 3445.550 ;
        RECT 1037.460 3435.000 1037.600 3445.230 ;
        RECT 1037.430 3431.000 1037.710 3435.000 ;
        RECT 2880.680 2435.750 2880.820 3445.230 ;
        RECT 2880.620 2435.430 2880.880 2435.750 ;
        RECT 2898.560 2435.430 2898.820 2435.750 ;
        RECT 2898.620 2434.245 2898.760 2435.430 ;
        RECT 2898.550 2433.875 2898.830 2434.245 ;
      LAYER via2 ;
        RECT 2898.550 2433.920 2898.830 2434.200 ;
      LAYER met3 ;
        RECT 2898.525 2434.210 2898.855 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2898.525 2433.910 2924.800 2434.210 ;
        RECT 2898.525 2433.895 2898.855 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 263.650 34.240 263.970 34.300 ;
        RECT 2902.670 34.240 2902.990 34.300 ;
        RECT 263.650 34.100 2902.990 34.240 ;
        RECT 263.650 34.040 263.970 34.100 ;
        RECT 2902.670 34.040 2902.990 34.100 ;
      LAYER via ;
        RECT 263.680 34.040 263.940 34.300 ;
        RECT 2902.700 34.040 2902.960 34.300 ;
      LAYER met2 ;
        RECT 2902.690 2669.155 2902.970 2669.525 ;
        RECT 263.710 35.000 263.990 39.000 ;
        RECT 263.740 34.330 263.880 35.000 ;
        RECT 2902.760 34.330 2902.900 2669.155 ;
        RECT 263.680 34.010 263.940 34.330 ;
        RECT 2902.700 34.010 2902.960 34.330 ;
      LAYER via2 ;
        RECT 2902.690 2669.200 2902.970 2669.480 ;
      LAYER met3 ;
        RECT 2902.665 2669.490 2902.995 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2902.665 2669.190 2924.800 2669.490 ;
        RECT 2902.665 2669.175 2902.995 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 314.710 33.900 315.030 33.960 ;
        RECT 2902.210 33.900 2902.530 33.960 ;
        RECT 314.710 33.760 2902.530 33.900 ;
        RECT 314.710 33.700 315.030 33.760 ;
        RECT 2902.210 33.700 2902.530 33.760 ;
      LAYER via ;
        RECT 314.740 33.700 315.000 33.960 ;
        RECT 2902.240 33.700 2902.500 33.960 ;
      LAYER met2 ;
        RECT 2902.230 2903.755 2902.510 2904.125 ;
        RECT 314.770 35.000 315.050 39.000 ;
        RECT 314.800 33.990 314.940 35.000 ;
        RECT 2902.300 33.990 2902.440 2903.755 ;
        RECT 314.740 33.670 315.000 33.990 ;
        RECT 2902.240 33.670 2902.500 33.990 ;
      LAYER via2 ;
        RECT 2902.230 2903.800 2902.510 2904.080 ;
      LAYER met3 ;
        RECT 2902.205 2904.090 2902.535 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2902.205 2903.790 2924.800 2904.090 ;
        RECT 2902.205 2903.775 2902.535 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 33.560 365.630 33.620 ;
        RECT 2901.750 33.560 2902.070 33.620 ;
        RECT 365.310 33.420 2902.070 33.560 ;
        RECT 365.310 33.360 365.630 33.420 ;
        RECT 2901.750 33.360 2902.070 33.420 ;
      LAYER via ;
        RECT 365.340 33.360 365.600 33.620 ;
        RECT 2901.780 33.360 2902.040 33.620 ;
      LAYER met2 ;
        RECT 2901.770 3138.355 2902.050 3138.725 ;
        RECT 365.370 35.000 365.650 39.000 ;
        RECT 365.400 33.650 365.540 35.000 ;
        RECT 2901.840 33.650 2901.980 3138.355 ;
        RECT 365.340 33.330 365.600 33.650 ;
        RECT 2901.780 33.330 2902.040 33.650 ;
      LAYER via2 ;
        RECT 2901.770 3138.400 2902.050 3138.680 ;
      LAYER met3 ;
        RECT 2901.745 3138.690 2902.075 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2901.745 3138.390 2924.800 3138.690 ;
        RECT 2901.745 3138.375 2902.075 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 416.370 33.220 416.690 33.280 ;
        RECT 2901.290 33.220 2901.610 33.280 ;
        RECT 416.370 33.080 2901.610 33.220 ;
        RECT 416.370 33.020 416.690 33.080 ;
        RECT 2901.290 33.020 2901.610 33.080 ;
      LAYER via ;
        RECT 416.400 33.020 416.660 33.280 ;
        RECT 2901.320 33.020 2901.580 33.280 ;
      LAYER met2 ;
        RECT 2901.310 3372.955 2901.590 3373.325 ;
        RECT 416.430 35.000 416.710 39.000 ;
        RECT 416.460 33.310 416.600 35.000 ;
        RECT 2901.380 33.310 2901.520 3372.955 ;
        RECT 416.400 32.990 416.660 33.310 ;
        RECT 2901.320 32.990 2901.580 33.310 ;
      LAYER via2 ;
        RECT 2901.310 3373.000 2901.590 3373.280 ;
      LAYER met3 ;
        RECT 2901.285 3373.290 2901.615 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2901.285 3372.990 2924.800 3373.290 ;
        RECT 2901.285 3372.975 2901.615 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 89.310 3501.560 89.630 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 89.310 3501.420 2798.570 3501.560 ;
        RECT 89.310 3501.360 89.630 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
      LAYER via ;
        RECT 89.340 3501.360 89.600 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 89.340 3501.330 89.600 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 87.530 3434.410 87.810 3435.000 ;
        RECT 89.400 3434.410 89.540 3501.330 ;
        RECT 87.530 3434.270 89.540 3434.410 ;
        RECT 87.530 3431.000 87.810 3434.270 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.810 3501.900 193.130 3501.960 ;
        RECT 2473.950 3501.900 2474.270 3501.960 ;
        RECT 192.810 3501.760 2474.270 3501.900 ;
        RECT 192.810 3501.700 193.130 3501.760 ;
        RECT 2473.950 3501.700 2474.270 3501.760 ;
      LAYER via ;
        RECT 192.840 3501.700 193.100 3501.960 ;
        RECT 2473.980 3501.700 2474.240 3501.960 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3501.990 2474.180 3517.600 ;
        RECT 192.840 3501.670 193.100 3501.990 ;
        RECT 2473.980 3501.670 2474.240 3501.990 ;
        RECT 192.900 3435.000 193.040 3501.670 ;
        RECT 192.870 3431.000 193.150 3435.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 303.210 3502.240 303.530 3502.300 ;
        RECT 2149.190 3502.240 2149.510 3502.300 ;
        RECT 303.210 3502.100 2149.510 3502.240 ;
        RECT 303.210 3502.040 303.530 3502.100 ;
        RECT 2149.190 3502.040 2149.510 3502.100 ;
        RECT 298.150 3448.520 298.470 3448.580 ;
        RECT 303.210 3448.520 303.530 3448.580 ;
        RECT 298.150 3448.380 303.530 3448.520 ;
        RECT 298.150 3448.320 298.470 3448.380 ;
        RECT 303.210 3448.320 303.530 3448.380 ;
      LAYER via ;
        RECT 303.240 3502.040 303.500 3502.300 ;
        RECT 2149.220 3502.040 2149.480 3502.300 ;
        RECT 298.180 3448.320 298.440 3448.580 ;
        RECT 303.240 3448.320 303.500 3448.580 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3502.330 2149.420 3517.600 ;
        RECT 303.240 3502.010 303.500 3502.330 ;
        RECT 2149.220 3502.010 2149.480 3502.330 ;
        RECT 303.300 3448.610 303.440 3502.010 ;
        RECT 298.180 3448.290 298.440 3448.610 ;
        RECT 303.240 3448.290 303.500 3448.610 ;
        RECT 298.240 3435.000 298.380 3448.290 ;
        RECT 298.210 3431.000 298.490 3435.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 406.710 3502.580 407.030 3502.640 ;
        RECT 1824.890 3502.580 1825.210 3502.640 ;
        RECT 406.710 3502.440 1825.210 3502.580 ;
        RECT 406.710 3502.380 407.030 3502.440 ;
        RECT 1824.890 3502.380 1825.210 3502.440 ;
      LAYER via ;
        RECT 406.740 3502.380 407.000 3502.640 ;
        RECT 1824.920 3502.380 1825.180 3502.640 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3502.670 1825.120 3517.600 ;
        RECT 406.740 3502.350 407.000 3502.670 ;
        RECT 1824.920 3502.350 1825.180 3502.670 ;
        RECT 404.010 3433.730 404.290 3435.000 ;
        RECT 406.800 3433.730 406.940 3502.350 ;
        RECT 404.010 3433.590 406.940 3433.730 ;
        RECT 404.010 3431.000 404.290 3433.590 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 510.210 3502.920 510.530 3502.980 ;
        RECT 1500.590 3502.920 1500.910 3502.980 ;
        RECT 510.210 3502.780 1500.910 3502.920 ;
        RECT 510.210 3502.720 510.530 3502.780 ;
        RECT 1500.590 3502.720 1500.910 3502.780 ;
      LAYER via ;
        RECT 510.240 3502.720 510.500 3502.980 ;
        RECT 1500.620 3502.720 1500.880 3502.980 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3503.010 1500.820 3517.600 ;
        RECT 510.240 3502.690 510.500 3503.010 ;
        RECT 1500.620 3502.690 1500.880 3503.010 ;
        RECT 509.350 3434.410 509.630 3435.000 ;
        RECT 510.300 3434.410 510.440 3502.690 ;
        RECT 509.350 3434.270 510.440 3434.410 ;
        RECT 509.350 3431.000 509.630 3434.270 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 220.220 2891.030 220.280 ;
        RECT 2903.130 220.220 2903.450 220.280 ;
        RECT 2890.710 220.080 2903.450 220.220 ;
        RECT 2890.710 220.020 2891.030 220.080 ;
        RECT 2903.130 220.020 2903.450 220.080 ;
      LAYER via ;
        RECT 2890.740 220.020 2891.000 220.280 ;
        RECT 2903.160 220.020 2903.420 220.280 ;
      LAYER met2 ;
        RECT 2903.150 322.475 2903.430 322.845 ;
        RECT 2903.220 220.310 2903.360 322.475 ;
        RECT 2890.740 220.165 2891.000 220.310 ;
        RECT 2890.730 219.795 2891.010 220.165 ;
        RECT 2903.160 219.990 2903.420 220.310 ;
      LAYER via2 ;
        RECT 2903.150 322.520 2903.430 322.800 ;
        RECT 2890.730 219.840 2891.010 220.120 ;
      LAYER met3 ;
        RECT 2903.125 322.810 2903.455 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2903.125 322.510 2924.800 322.810 ;
        RECT 2903.125 322.495 2903.455 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
        RECT 2890.705 220.130 2891.035 220.145 ;
        RECT 2884.510 219.830 2891.035 220.130 ;
        RECT 2884.510 217.200 2884.810 219.830 ;
        RECT 2890.705 219.815 2891.035 219.830 ;
        RECT 2881.000 216.600 2885.000 217.200 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 620.610 3503.260 620.930 3503.320 ;
        RECT 1175.830 3503.260 1176.150 3503.320 ;
        RECT 620.610 3503.120 1176.150 3503.260 ;
        RECT 620.610 3503.060 620.930 3503.120 ;
        RECT 1175.830 3503.060 1176.150 3503.120 ;
        RECT 615.090 3448.860 615.410 3448.920 ;
        RECT 620.610 3448.860 620.930 3448.920 ;
        RECT 615.090 3448.720 620.930 3448.860 ;
        RECT 615.090 3448.660 615.410 3448.720 ;
        RECT 620.610 3448.660 620.930 3448.720 ;
      LAYER via ;
        RECT 620.640 3503.060 620.900 3503.320 ;
        RECT 1175.860 3503.060 1176.120 3503.320 ;
        RECT 615.120 3448.660 615.380 3448.920 ;
        RECT 620.640 3448.660 620.900 3448.920 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3503.350 1176.060 3517.600 ;
        RECT 620.640 3503.030 620.900 3503.350 ;
        RECT 1175.860 3503.030 1176.120 3503.350 ;
        RECT 620.700 3448.950 620.840 3503.030 ;
        RECT 615.120 3448.630 615.380 3448.950 ;
        RECT 620.640 3448.630 620.900 3448.950 ;
        RECT 615.180 3435.000 615.320 3448.630 ;
        RECT 615.150 3431.000 615.430 3435.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 724.110 3503.600 724.430 3503.660 ;
        RECT 851.530 3503.600 851.850 3503.660 ;
        RECT 724.110 3503.460 851.850 3503.600 ;
        RECT 724.110 3503.400 724.430 3503.460 ;
        RECT 851.530 3503.400 851.850 3503.460 ;
        RECT 720.430 3448.860 720.750 3448.920 ;
        RECT 724.110 3448.860 724.430 3448.920 ;
        RECT 720.430 3448.720 724.430 3448.860 ;
        RECT 720.430 3448.660 720.750 3448.720 ;
        RECT 724.110 3448.660 724.430 3448.720 ;
      LAYER via ;
        RECT 724.140 3503.400 724.400 3503.660 ;
        RECT 851.560 3503.400 851.820 3503.660 ;
        RECT 720.460 3448.660 720.720 3448.920 ;
        RECT 724.140 3448.660 724.400 3448.920 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3503.690 851.760 3517.600 ;
        RECT 724.140 3503.370 724.400 3503.690 ;
        RECT 851.560 3503.370 851.820 3503.690 ;
        RECT 724.200 3448.950 724.340 3503.370 ;
        RECT 720.460 3448.630 720.720 3448.950 ;
        RECT 724.140 3448.630 724.400 3448.950 ;
        RECT 720.520 3435.000 720.660 3448.630 ;
        RECT 720.490 3431.000 720.770 3435.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3503.260 527.550 3503.320 ;
        RECT 530.910 3503.260 531.230 3503.320 ;
        RECT 527.230 3503.120 531.230 3503.260 ;
        RECT 527.230 3503.060 527.550 3503.120 ;
        RECT 530.910 3503.060 531.230 3503.120 ;
        RECT 530.910 3448.520 531.230 3448.580 ;
        RECT 826.230 3448.520 826.550 3448.580 ;
        RECT 530.910 3448.380 826.550 3448.520 ;
        RECT 530.910 3448.320 531.230 3448.380 ;
        RECT 826.230 3448.320 826.550 3448.380 ;
      LAYER via ;
        RECT 527.260 3503.060 527.520 3503.320 ;
        RECT 530.940 3503.060 531.200 3503.320 ;
        RECT 530.940 3448.320 531.200 3448.580 ;
        RECT 826.260 3448.320 826.520 3448.580 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.350 527.460 3517.600 ;
        RECT 527.260 3503.030 527.520 3503.350 ;
        RECT 530.940 3503.030 531.200 3503.350 ;
        RECT 531.000 3448.610 531.140 3503.030 ;
        RECT 530.940 3448.290 531.200 3448.610 ;
        RECT 826.260 3448.290 826.520 3448.610 ;
        RECT 826.320 3435.000 826.460 3448.290 ;
        RECT 826.290 3431.000 826.570 3435.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.240 202.790 3502.300 ;
        RECT 206.610 3502.240 206.930 3502.300 ;
        RECT 202.470 3502.100 206.930 3502.240 ;
        RECT 202.470 3502.040 202.790 3502.100 ;
        RECT 206.610 3502.040 206.930 3502.100 ;
        RECT 206.610 3448.180 206.930 3448.240 ;
        RECT 931.570 3448.180 931.890 3448.240 ;
        RECT 206.610 3448.040 931.890 3448.180 ;
        RECT 206.610 3447.980 206.930 3448.040 ;
        RECT 931.570 3447.980 931.890 3448.040 ;
      LAYER via ;
        RECT 202.500 3502.040 202.760 3502.300 ;
        RECT 206.640 3502.040 206.900 3502.300 ;
        RECT 206.640 3447.980 206.900 3448.240 ;
        RECT 931.600 3447.980 931.860 3448.240 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3502.330 202.700 3517.600 ;
        RECT 202.500 3502.010 202.760 3502.330 ;
        RECT 206.640 3502.010 206.900 3502.330 ;
        RECT 206.700 3448.270 206.840 3502.010 ;
        RECT 206.640 3447.950 206.900 3448.270 ;
        RECT 931.600 3447.950 931.860 3448.270 ;
        RECT 931.660 3435.000 931.800 3447.950 ;
        RECT 931.630 3431.000 931.910 3435.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.710 3408.740 16.030 3408.800 ;
        RECT 30.890 3408.740 31.210 3408.800 ;
        RECT 15.710 3408.600 31.210 3408.740 ;
        RECT 15.710 3408.540 16.030 3408.600 ;
        RECT 30.890 3408.540 31.210 3408.600 ;
        RECT 30.890 26.420 31.210 26.480 ;
        RECT 60.330 26.420 60.650 26.480 ;
        RECT 30.890 26.280 60.650 26.420 ;
        RECT 30.890 26.220 31.210 26.280 ;
        RECT 60.330 26.220 60.650 26.280 ;
      LAYER via ;
        RECT 15.740 3408.540 16.000 3408.800 ;
        RECT 30.920 3408.540 31.180 3408.800 ;
        RECT 30.920 26.220 31.180 26.480 ;
        RECT 60.360 26.220 60.620 26.480 ;
      LAYER met2 ;
        RECT 15.730 3411.035 16.010 3411.405 ;
        RECT 15.800 3408.830 15.940 3411.035 ;
        RECT 15.740 3408.510 16.000 3408.830 ;
        RECT 30.920 3408.510 31.180 3408.830 ;
        RECT 30.980 26.510 31.120 3408.510 ;
        RECT 60.390 35.000 60.670 39.000 ;
        RECT 60.420 26.510 60.560 35.000 ;
        RECT 30.920 26.190 31.180 26.510 ;
        RECT 60.360 26.190 60.620 26.510 ;
      LAYER via2 ;
        RECT 15.730 3411.080 16.010 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 15.705 3411.370 16.035 3411.385 ;
        RECT -4.800 3411.070 16.035 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 15.705 3411.055 16.035 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 26.760 17.410 26.820 ;
        RECT 110.930 26.760 111.250 26.820 ;
        RECT 17.090 26.620 111.250 26.760 ;
        RECT 17.090 26.560 17.410 26.620 ;
        RECT 110.930 26.560 111.250 26.620 ;
      LAYER via ;
        RECT 17.120 26.560 17.380 26.820 ;
        RECT 110.960 26.560 111.220 26.820 ;
      LAYER met2 ;
        RECT 17.110 3124.075 17.390 3124.445 ;
        RECT 17.180 26.850 17.320 3124.075 ;
        RECT 110.990 35.000 111.270 39.000 ;
        RECT 111.020 26.850 111.160 35.000 ;
        RECT 17.120 26.530 17.380 26.850 ;
        RECT 110.960 26.530 111.220 26.850 ;
      LAYER via2 ;
        RECT 17.110 3124.120 17.390 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.085 3124.410 17.415 3124.425 ;
        RECT -4.800 3124.110 17.415 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.085 3124.095 17.415 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.850 2836.180 20.170 2836.240 ;
        RECT 31.350 2836.180 31.670 2836.240 ;
        RECT 19.850 2836.040 31.670 2836.180 ;
        RECT 19.850 2835.980 20.170 2836.040 ;
        RECT 31.350 2835.980 31.670 2836.040 ;
        RECT 31.350 27.100 31.670 27.160 ;
        RECT 161.990 27.100 162.310 27.160 ;
        RECT 31.350 26.960 162.310 27.100 ;
        RECT 31.350 26.900 31.670 26.960 ;
        RECT 161.990 26.900 162.310 26.960 ;
      LAYER via ;
        RECT 19.880 2835.980 20.140 2836.240 ;
        RECT 31.380 2835.980 31.640 2836.240 ;
        RECT 31.380 26.900 31.640 27.160 ;
        RECT 162.020 26.900 162.280 27.160 ;
      LAYER met2 ;
        RECT 19.870 2836.435 20.150 2836.805 ;
        RECT 19.940 2836.270 20.080 2836.435 ;
        RECT 19.880 2835.950 20.140 2836.270 ;
        RECT 31.380 2835.950 31.640 2836.270 ;
        RECT 31.440 27.190 31.580 2835.950 ;
        RECT 162.050 35.000 162.330 39.000 ;
        RECT 162.080 27.190 162.220 35.000 ;
        RECT 31.380 26.870 31.640 27.190 ;
        RECT 162.020 26.870 162.280 27.190 ;
      LAYER via2 ;
        RECT 19.870 2836.480 20.150 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 19.845 2836.770 20.175 2836.785 ;
        RECT -4.800 2836.470 20.175 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 19.845 2836.455 20.175 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 2546.500 17.870 2546.560 ;
        RECT 37.790 2546.500 38.110 2546.560 ;
        RECT 17.550 2546.360 38.110 2546.500 ;
        RECT 17.550 2546.300 17.870 2546.360 ;
        RECT 37.790 2546.300 38.110 2546.360 ;
        RECT 37.790 27.440 38.110 27.500 ;
        RECT 212.590 27.440 212.910 27.500 ;
        RECT 37.790 27.300 212.910 27.440 ;
        RECT 37.790 27.240 38.110 27.300 ;
        RECT 212.590 27.240 212.910 27.300 ;
      LAYER via ;
        RECT 17.580 2546.300 17.840 2546.560 ;
        RECT 37.820 2546.300 38.080 2546.560 ;
        RECT 37.820 27.240 38.080 27.500 ;
        RECT 212.620 27.240 212.880 27.500 ;
      LAYER met2 ;
        RECT 17.570 2549.475 17.850 2549.845 ;
        RECT 17.640 2546.590 17.780 2549.475 ;
        RECT 17.580 2546.270 17.840 2546.590 ;
        RECT 37.820 2546.270 38.080 2546.590 ;
        RECT 37.880 27.530 38.020 2546.270 ;
        RECT 212.650 35.000 212.930 39.000 ;
        RECT 212.680 27.530 212.820 35.000 ;
        RECT 37.820 27.210 38.080 27.530 ;
        RECT 212.620 27.210 212.880 27.530 ;
      LAYER via2 ;
        RECT 17.570 2549.520 17.850 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 17.545 2549.810 17.875 2549.825 ;
        RECT -4.800 2549.510 17.875 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 17.545 2549.495 17.875 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 2261.835 17.850 2262.205 ;
        RECT 17.640 89.605 17.780 2261.835 ;
        RECT 17.570 89.235 17.850 89.605 ;
      LAYER via2 ;
        RECT 17.570 2261.880 17.850 2262.160 ;
        RECT 17.570 89.280 17.850 89.560 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.545 2262.170 17.875 2262.185 ;
        RECT -4.800 2261.870 17.875 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.545 2261.855 17.875 2261.870 ;
        RECT 17.545 89.570 17.875 89.585 ;
        RECT 17.545 89.270 35.570 89.570 ;
        RECT 17.545 89.255 17.875 89.270 ;
        RECT 35.270 86.640 35.570 89.270 ;
        RECT 35.000 86.040 39.000 86.640 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 1974.875 18.310 1975.245 ;
        RECT 18.100 191.605 18.240 1974.875 ;
        RECT 18.030 191.235 18.310 191.605 ;
      LAYER via2 ;
        RECT 18.030 1974.920 18.310 1975.200 ;
        RECT 18.030 191.280 18.310 191.560 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 18.005 1975.210 18.335 1975.225 ;
        RECT -4.800 1974.910 18.335 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 18.005 1974.895 18.335 1974.910 ;
        RECT 18.005 191.570 18.335 191.585 ;
        RECT 18.005 191.270 35.570 191.570 ;
        RECT 18.005 191.255 18.335 191.270 ;
        RECT 35.270 189.320 35.570 191.270 ;
        RECT 35.000 188.720 39.000 189.320 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 341.940 2891.030 342.000 ;
        RECT 2903.130 341.940 2903.450 342.000 ;
        RECT 2890.710 341.800 2903.450 341.940 ;
        RECT 2890.710 341.740 2891.030 341.800 ;
        RECT 2903.130 341.740 2903.450 341.800 ;
      LAYER via ;
        RECT 2890.740 341.740 2891.000 342.000 ;
        RECT 2903.160 341.740 2903.420 342.000 ;
      LAYER met2 ;
        RECT 2903.150 557.075 2903.430 557.445 ;
        RECT 2903.220 342.030 2903.360 557.075 ;
        RECT 2890.740 341.885 2891.000 342.030 ;
        RECT 2890.730 341.515 2891.010 341.885 ;
        RECT 2903.160 341.710 2903.420 342.030 ;
      LAYER via2 ;
        RECT 2903.150 557.120 2903.430 557.400 ;
        RECT 2890.730 341.560 2891.010 341.840 ;
      LAYER met3 ;
        RECT 2903.125 557.410 2903.455 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2903.125 557.110 2924.800 557.410 ;
        RECT 2903.125 557.095 2903.455 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
        RECT 2890.705 341.850 2891.035 341.865 ;
        RECT 2884.510 341.550 2891.035 341.850 ;
        RECT 2884.510 338.920 2884.810 341.550 ;
        RECT 2890.705 341.535 2891.035 341.550 ;
        RECT 2881.000 338.320 2885.000 338.920 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 1687.235 18.770 1687.605 ;
        RECT 18.560 295.645 18.700 1687.235 ;
        RECT 18.490 295.275 18.770 295.645 ;
      LAYER via2 ;
        RECT 18.490 1687.280 18.770 1687.560 ;
        RECT 18.490 295.320 18.770 295.600 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 18.465 1687.570 18.795 1687.585 ;
        RECT -4.800 1687.270 18.795 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 18.465 1687.255 18.795 1687.270 ;
        RECT 18.465 295.610 18.795 295.625 ;
        RECT 18.465 295.310 35.570 295.610 ;
        RECT 18.465 295.295 18.795 295.310 ;
        RECT 35.270 292.680 35.570 295.310 ;
        RECT 35.000 292.080 39.000 292.680 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 1471.675 19.230 1472.045 ;
        RECT 19.020 398.325 19.160 1471.675 ;
        RECT 18.950 397.955 19.230 398.325 ;
      LAYER via2 ;
        RECT 18.950 1471.720 19.230 1472.000 ;
        RECT 18.950 398.000 19.230 398.280 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 18.925 1472.010 19.255 1472.025 ;
        RECT -4.800 1471.710 19.255 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 18.925 1471.695 19.255 1471.710 ;
        RECT 18.925 398.290 19.255 398.305 ;
        RECT 18.925 397.990 35.570 398.290 ;
        RECT 18.925 397.975 19.255 397.990 ;
        RECT 35.270 395.360 35.570 397.990 ;
        RECT 35.000 394.760 39.000 395.360 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 1256.115 20.150 1256.485 ;
        RECT 19.940 501.685 20.080 1256.115 ;
        RECT 19.870 501.315 20.150 501.685 ;
      LAYER via2 ;
        RECT 19.870 1256.160 20.150 1256.440 ;
        RECT 19.870 501.360 20.150 501.640 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 19.845 1256.450 20.175 1256.465 ;
        RECT -4.800 1256.150 20.175 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 19.845 1256.135 20.175 1256.150 ;
        RECT 19.845 501.650 20.175 501.665 ;
        RECT 19.845 501.350 35.570 501.650 ;
        RECT 19.845 501.335 20.175 501.350 ;
        RECT 35.270 498.720 35.570 501.350 ;
        RECT 35.000 498.120 39.000 498.720 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 607.140 16.490 607.200 ;
        RECT 20.770 607.140 21.090 607.200 ;
        RECT 16.170 607.000 21.090 607.140 ;
        RECT 16.170 606.940 16.490 607.000 ;
        RECT 20.770 606.940 21.090 607.000 ;
      LAYER via ;
        RECT 16.200 606.940 16.460 607.200 ;
        RECT 20.800 606.940 21.060 607.200 ;
      LAYER met2 ;
        RECT 16.190 1040.555 16.470 1040.925 ;
        RECT 16.260 607.230 16.400 1040.555 ;
        RECT 16.200 606.910 16.460 607.230 ;
        RECT 20.800 606.910 21.060 607.230 ;
        RECT 20.860 604.365 21.000 606.910 ;
        RECT 20.790 603.995 21.070 604.365 ;
      LAYER via2 ;
        RECT 16.190 1040.600 16.470 1040.880 ;
        RECT 20.790 604.040 21.070 604.320 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 16.165 1040.890 16.495 1040.905 ;
        RECT -4.800 1040.590 16.495 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 16.165 1040.575 16.495 1040.590 ;
        RECT 20.765 604.330 21.095 604.345 ;
        RECT 20.765 604.030 35.570 604.330 ;
        RECT 20.765 604.015 21.095 604.030 ;
        RECT 35.270 601.400 35.570 604.030 ;
        RECT 35.000 600.800 39.000 601.400 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.730 824.995 16.010 825.365 ;
        RECT 15.800 707.725 15.940 824.995 ;
        RECT 15.730 707.355 16.010 707.725 ;
      LAYER via2 ;
        RECT 15.730 825.040 16.010 825.320 ;
        RECT 15.730 707.400 16.010 707.680 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 15.705 825.330 16.035 825.345 ;
        RECT -4.800 825.030 16.035 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 15.705 825.015 16.035 825.030 ;
        RECT 15.705 707.690 16.035 707.705 ;
        RECT 15.705 707.390 35.570 707.690 ;
        RECT 15.705 707.375 16.035 707.390 ;
        RECT 35.270 704.760 35.570 707.390 ;
        RECT 35.000 704.160 39.000 704.760 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 803.915 21.070 804.285 ;
        RECT 20.860 610.485 21.000 803.915 ;
        RECT 20.790 610.115 21.070 610.485 ;
      LAYER via2 ;
        RECT 20.790 803.960 21.070 804.240 ;
        RECT 20.790 610.160 21.070 610.440 ;
      LAYER met3 ;
        RECT 35.000 806.840 39.000 807.440 ;
        RECT 20.765 804.250 21.095 804.265 ;
        RECT 35.270 804.250 35.570 806.840 ;
        RECT 20.765 803.950 35.570 804.250 ;
        RECT 20.765 803.935 21.095 803.950 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 20.765 610.450 21.095 610.465 ;
        RECT -4.800 610.150 21.095 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 20.765 610.135 21.095 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 905.660 16.950 905.720 ;
        RECT 20.770 905.660 21.090 905.720 ;
        RECT 16.630 905.520 21.090 905.660 ;
        RECT 16.630 905.460 16.950 905.520 ;
        RECT 20.770 905.460 21.090 905.520 ;
      LAYER via ;
        RECT 16.660 905.460 16.920 905.720 ;
        RECT 20.800 905.460 21.060 905.720 ;
      LAYER met2 ;
        RECT 20.790 907.275 21.070 907.645 ;
        RECT 20.860 905.750 21.000 907.275 ;
        RECT 16.660 905.430 16.920 905.750 ;
        RECT 20.800 905.430 21.060 905.750 ;
        RECT 16.720 394.925 16.860 905.430 ;
        RECT 16.650 394.555 16.930 394.925 ;
      LAYER via2 ;
        RECT 20.790 907.320 21.070 907.600 ;
        RECT 16.650 394.600 16.930 394.880 ;
      LAYER met3 ;
        RECT 35.000 910.200 39.000 910.800 ;
        RECT 20.765 907.610 21.095 907.625 ;
        RECT 35.270 907.610 35.570 910.200 ;
        RECT 20.765 907.310 35.570 907.610 ;
        RECT 20.765 907.295 21.095 907.310 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 16.625 394.890 16.955 394.905 ;
        RECT -4.800 394.590 16.955 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 16.625 394.575 16.955 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 1009.955 19.690 1010.325 ;
        RECT 19.480 179.365 19.620 1009.955 ;
        RECT 19.410 178.995 19.690 179.365 ;
      LAYER via2 ;
        RECT 19.410 1010.000 19.690 1010.280 ;
        RECT 19.410 179.040 19.690 179.320 ;
      LAYER met3 ;
        RECT 35.000 1012.880 39.000 1013.480 ;
        RECT 19.385 1010.290 19.715 1010.305 ;
        RECT 35.270 1010.290 35.570 1012.880 ;
        RECT 19.385 1009.990 35.570 1010.290 ;
        RECT 19.385 1009.975 19.715 1009.990 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 19.385 179.330 19.715 179.345 ;
        RECT -4.800 179.030 19.715 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 19.385 179.015 19.715 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 462.300 2891.030 462.360 ;
        RECT 2903.590 462.300 2903.910 462.360 ;
        RECT 2890.710 462.160 2903.910 462.300 ;
        RECT 2890.710 462.100 2891.030 462.160 ;
        RECT 2903.590 462.100 2903.910 462.160 ;
      LAYER via ;
        RECT 2890.740 462.100 2891.000 462.360 ;
        RECT 2903.620 462.100 2903.880 462.360 ;
      LAYER met2 ;
        RECT 2903.610 791.675 2903.890 792.045 ;
        RECT 2903.680 462.390 2903.820 791.675 ;
        RECT 2890.740 462.245 2891.000 462.390 ;
        RECT 2890.730 461.875 2891.010 462.245 ;
        RECT 2903.620 462.070 2903.880 462.390 ;
      LAYER via2 ;
        RECT 2903.610 791.720 2903.890 792.000 ;
        RECT 2890.730 461.920 2891.010 462.200 ;
      LAYER met3 ;
        RECT 2903.585 792.010 2903.915 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2903.585 791.710 2924.800 792.010 ;
        RECT 2903.585 791.695 2903.915 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
        RECT 2890.705 462.210 2891.035 462.225 ;
        RECT 2884.510 461.910 2891.035 462.210 ;
        RECT 2884.510 459.960 2884.810 461.910 ;
        RECT 2890.705 461.895 2891.035 461.910 ;
        RECT 2881.000 459.360 2885.000 459.960 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 584.700 2891.030 584.760 ;
        RECT 2903.130 584.700 2903.450 584.760 ;
        RECT 2890.710 584.560 2903.450 584.700 ;
        RECT 2890.710 584.500 2891.030 584.560 ;
        RECT 2903.130 584.500 2903.450 584.560 ;
      LAYER via ;
        RECT 2890.740 584.500 2891.000 584.760 ;
        RECT 2903.160 584.500 2903.420 584.760 ;
      LAYER met2 ;
        RECT 2903.150 1026.275 2903.430 1026.645 ;
        RECT 2903.220 584.790 2903.360 1026.275 ;
        RECT 2890.740 584.645 2891.000 584.790 ;
        RECT 2890.730 584.275 2891.010 584.645 ;
        RECT 2903.160 584.470 2903.420 584.790 ;
      LAYER via2 ;
        RECT 2903.150 1026.320 2903.430 1026.600 ;
        RECT 2890.730 584.320 2891.010 584.600 ;
      LAYER met3 ;
        RECT 2903.125 1026.610 2903.455 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2903.125 1026.310 2924.800 1026.610 ;
        RECT 2903.125 1026.295 2903.455 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
        RECT 2890.705 584.610 2891.035 584.625 ;
        RECT 2884.510 584.310 2891.035 584.610 ;
        RECT 2884.510 581.680 2884.810 584.310 ;
        RECT 2890.705 584.295 2891.035 584.310 ;
        RECT 2881.000 581.080 2885.000 581.680 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2900.850 1260.875 2901.130 1261.245 ;
        RECT 2900.920 703.645 2901.060 1260.875 ;
        RECT 2900.850 703.275 2901.130 703.645 ;
      LAYER via2 ;
        RECT 2900.850 1260.920 2901.130 1261.200 ;
        RECT 2900.850 703.320 2901.130 703.600 ;
      LAYER met3 ;
        RECT 2900.825 1261.210 2901.155 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2900.825 1260.910 2924.800 1261.210 ;
        RECT 2900.825 1260.895 2901.155 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 2900.825 703.610 2901.155 703.625 ;
        RECT 2884.510 703.310 2901.155 703.610 ;
        RECT 2884.510 702.720 2884.810 703.310 ;
        RECT 2900.825 703.295 2901.155 703.310 ;
        RECT 2881.000 702.120 2885.000 702.720 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 827.460 2891.030 827.520 ;
        RECT 2904.510 827.460 2904.830 827.520 ;
        RECT 2890.710 827.320 2904.830 827.460 ;
        RECT 2890.710 827.260 2891.030 827.320 ;
        RECT 2904.510 827.260 2904.830 827.320 ;
      LAYER via ;
        RECT 2890.740 827.260 2891.000 827.520 ;
        RECT 2904.540 827.260 2904.800 827.520 ;
      LAYER met2 ;
        RECT 2904.530 1495.475 2904.810 1495.845 ;
        RECT 2904.600 827.550 2904.740 1495.475 ;
        RECT 2890.740 827.405 2891.000 827.550 ;
        RECT 2890.730 827.035 2891.010 827.405 ;
        RECT 2904.540 827.230 2904.800 827.550 ;
      LAYER via2 ;
        RECT 2904.530 1495.520 2904.810 1495.800 ;
        RECT 2890.730 827.080 2891.010 827.360 ;
      LAYER met3 ;
        RECT 2904.505 1495.810 2904.835 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2904.505 1495.510 2924.800 1495.810 ;
        RECT 2904.505 1495.495 2904.835 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2890.705 827.370 2891.035 827.385 ;
        RECT 2884.510 827.070 2891.035 827.370 ;
        RECT 2884.510 824.440 2884.810 827.070 ;
        RECT 2890.705 827.055 2891.035 827.070 ;
        RECT 2881.000 823.840 2885.000 824.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 949.180 2891.030 949.240 ;
        RECT 2904.050 949.180 2904.370 949.240 ;
        RECT 2890.710 949.040 2904.370 949.180 ;
        RECT 2890.710 948.980 2891.030 949.040 ;
        RECT 2904.050 948.980 2904.370 949.040 ;
      LAYER via ;
        RECT 2890.740 948.980 2891.000 949.240 ;
        RECT 2904.080 948.980 2904.340 949.240 ;
      LAYER met2 ;
        RECT 2904.070 1730.075 2904.350 1730.445 ;
        RECT 2904.140 949.270 2904.280 1730.075 ;
        RECT 2890.740 949.125 2891.000 949.270 ;
        RECT 2890.730 948.755 2891.010 949.125 ;
        RECT 2904.080 948.950 2904.340 949.270 ;
      LAYER via2 ;
        RECT 2904.070 1730.120 2904.350 1730.400 ;
        RECT 2890.730 948.800 2891.010 949.080 ;
      LAYER met3 ;
        RECT 2904.045 1730.410 2904.375 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2904.045 1730.110 2924.800 1730.410 ;
        RECT 2904.045 1730.095 2904.375 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2890.705 949.090 2891.035 949.105 ;
        RECT 2884.510 948.790 2891.035 949.090 ;
        RECT 2884.510 946.160 2884.810 948.790 ;
        RECT 2890.705 948.775 2891.035 948.790 ;
        RECT 2881.000 945.560 2885.000 946.160 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 1069.540 2891.030 1069.600 ;
        RECT 2903.590 1069.540 2903.910 1069.600 ;
        RECT 2890.710 1069.400 2903.910 1069.540 ;
        RECT 2890.710 1069.340 2891.030 1069.400 ;
        RECT 2903.590 1069.340 2903.910 1069.400 ;
      LAYER via ;
        RECT 2890.740 1069.340 2891.000 1069.600 ;
        RECT 2903.620 1069.340 2903.880 1069.600 ;
      LAYER met2 ;
        RECT 2903.610 1964.675 2903.890 1965.045 ;
        RECT 2903.680 1069.630 2903.820 1964.675 ;
        RECT 2890.740 1069.485 2891.000 1069.630 ;
        RECT 2890.730 1069.115 2891.010 1069.485 ;
        RECT 2903.620 1069.310 2903.880 1069.630 ;
      LAYER via2 ;
        RECT 2903.610 1964.720 2903.890 1965.000 ;
        RECT 2890.730 1069.160 2891.010 1069.440 ;
      LAYER met3 ;
        RECT 2903.585 1965.010 2903.915 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2903.585 1964.710 2924.800 1965.010 ;
        RECT 2903.585 1964.695 2903.915 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2890.705 1069.450 2891.035 1069.465 ;
        RECT 2884.510 1069.150 2891.035 1069.450 ;
        RECT 2884.510 1067.200 2884.810 1069.150 ;
        RECT 2890.705 1069.135 2891.035 1069.150 ;
        RECT 2881.000 1066.600 2885.000 1067.200 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2890.710 1191.260 2891.030 1191.320 ;
        RECT 2903.130 1191.260 2903.450 1191.320 ;
        RECT 2890.710 1191.120 2903.450 1191.260 ;
        RECT 2890.710 1191.060 2891.030 1191.120 ;
        RECT 2903.130 1191.060 2903.450 1191.120 ;
      LAYER via ;
        RECT 2890.740 1191.060 2891.000 1191.320 ;
        RECT 2903.160 1191.060 2903.420 1191.320 ;
      LAYER met2 ;
        RECT 2903.150 2199.275 2903.430 2199.645 ;
        RECT 2903.220 1191.350 2903.360 2199.275 ;
        RECT 2890.740 1191.205 2891.000 1191.350 ;
        RECT 2890.730 1190.835 2891.010 1191.205 ;
        RECT 2903.160 1191.030 2903.420 1191.350 ;
      LAYER via2 ;
        RECT 2903.150 2199.320 2903.430 2199.600 ;
        RECT 2890.730 1190.880 2891.010 1191.160 ;
      LAYER met3 ;
        RECT 2903.125 2199.610 2903.455 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2903.125 2199.310 2924.800 2199.610 ;
        RECT 2903.125 2199.295 2903.455 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2890.705 1191.170 2891.035 1191.185 ;
        RECT 2884.510 1190.870 2891.035 1191.170 ;
        RECT 2884.510 1188.920 2884.810 1190.870 ;
        RECT 2890.705 1190.855 2891.035 1190.870 ;
        RECT 2881.000 1188.320 2885.000 1188.920 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2551.100 2924.800 2552.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2785.700 2924.800 2786.900 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3254.900 2924.800 3256.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3489.500 2924.800 3490.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 2.400 3268.340 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2979.500 2.400 2980.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2692.540 2.400 2693.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2404.900 2.400 2406.100 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.940 2.400 2119.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 2.400 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 2.400 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 2.400 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 2.400 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 2.400 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 2.400 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 2.400 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 2.400 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 2.400 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2316.500 2924.800 2317.700 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2727.220 2924.800 2728.420 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2961.820 2924.800 2963.020 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3431.020 2924.800 3432.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3339.220 2.400 3340.420 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 3051.580 2.400 3052.780 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2764.620 2.400 2765.820 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2476.980 2.400 2478.180 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 2189.340 2.400 2190.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 2.400 1903.580 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1614.740 2.400 1615.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 1184.300 2.400 1185.500 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 2.400 969.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 753.180 2.400 754.380 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 537.620 2.400 538.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 322.060 2.400 323.260 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT -4.800 106.500 2.400 107.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2.830 24.040 3.150 24.100 ;
        RECT 2095.830 24.040 2096.150 24.100 ;
        RECT 2.830 23.900 2096.150 24.040 ;
        RECT 2.830 23.840 3.150 23.900 ;
        RECT 2095.830 23.840 2096.150 23.900 ;
      LAYER via ;
        RECT 2.860 23.840 3.120 24.100 ;
        RECT 2095.860 23.840 2096.120 24.100 ;
      LAYER met2 ;
        RECT 2095.890 35.000 2096.170 39.000 ;
        RECT 2095.920 24.130 2096.060 35.000 ;
        RECT 2.860 23.810 3.120 24.130 ;
        RECT 2095.860 23.810 2096.120 24.130 ;
        RECT 2.920 2.400 3.060 23.810 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 13.410 3447.840 13.730 3447.900 ;
        RECT 1142.710 3447.840 1143.030 3447.900 ;
        RECT 13.410 3447.700 1143.030 3447.840 ;
        RECT 13.410 3447.640 13.730 3447.700 ;
        RECT 1142.710 3447.640 1143.030 3447.700 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 13.410 17.580 13.730 17.640 ;
        RECT 8.350 17.440 13.730 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 13.410 17.380 13.730 17.440 ;
      LAYER via ;
        RECT 13.440 3447.640 13.700 3447.900 ;
        RECT 1142.740 3447.640 1143.000 3447.900 ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 13.440 17.380 13.700 17.640 ;
      LAYER met2 ;
        RECT 13.440 3447.610 13.700 3447.930 ;
        RECT 1142.740 3447.610 1143.000 3447.930 ;
        RECT 13.500 17.670 13.640 3447.610 ;
        RECT 1142.800 3435.000 1142.940 3447.610 ;
        RECT 1142.770 3431.000 1143.050 3435.000 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 13.440 17.350 13.700 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2146.950 35.000 2147.230 39.000 ;
        RECT 2146.980 27.045 2147.120 35.000 ;
        RECT 14.350 26.675 14.630 27.045 ;
        RECT 2146.910 26.675 2147.190 27.045 ;
        RECT 14.420 2.400 14.560 26.675 ;
        RECT 14.210 -4.800 14.770 2.400 ;
      LAYER via2 ;
        RECT 14.350 26.720 14.630 27.000 ;
        RECT 2146.910 26.720 2147.190 27.000 ;
      LAYER met3 ;
        RECT 14.325 27.010 14.655 27.025 ;
        RECT 2146.885 27.010 2147.215 27.025 ;
        RECT 14.325 26.710 2147.215 27.010 ;
        RECT 14.325 26.695 14.655 26.710 ;
        RECT 2146.885 26.695 2147.215 26.710 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.970 1113.315 36.250 1113.685 ;
        RECT 36.040 16.050 36.180 1113.315 ;
        RECT 36.040 15.910 38.480 16.050 ;
        RECT 38.340 2.400 38.480 15.910 ;
        RECT 38.130 -4.800 38.690 2.400 ;
      LAYER via2 ;
        RECT 35.970 1113.360 36.250 1113.640 ;
      LAYER met3 ;
        RECT 35.000 1116.240 39.000 1116.840 ;
        RECT 36.190 1113.665 36.490 1116.240 ;
        RECT 35.945 1113.350 36.490 1113.665 ;
        RECT 35.945 1113.335 36.275 1113.350 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 240.650 25.060 240.970 25.120 ;
        RECT 2248.550 25.060 2248.870 25.120 ;
        RECT 240.650 24.920 2248.870 25.060 ;
        RECT 240.650 24.860 240.970 24.920 ;
        RECT 2248.550 24.860 2248.870 24.920 ;
      LAYER via ;
        RECT 240.680 24.860 240.940 25.120 ;
        RECT 2248.580 24.860 2248.840 25.120 ;
      LAYER met2 ;
        RECT 2248.610 35.000 2248.890 39.000 ;
        RECT 2248.640 25.150 2248.780 35.000 ;
        RECT 240.680 24.830 240.940 25.150 ;
        RECT 2248.580 24.830 2248.840 25.150 ;
        RECT 240.740 2.400 240.880 24.830 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 21.230 24.720 21.550 24.780 ;
        RECT 258.130 24.720 258.450 24.780 ;
        RECT 21.230 24.580 258.450 24.720 ;
        RECT 21.230 24.520 21.550 24.580 ;
        RECT 258.130 24.520 258.450 24.580 ;
      LAYER via ;
        RECT 21.260 24.520 21.520 24.780 ;
        RECT 258.160 24.520 258.420 24.780 ;
      LAYER met2 ;
        RECT 21.250 1628.755 21.530 1629.125 ;
        RECT 21.320 24.810 21.460 1628.755 ;
        RECT 21.260 24.490 21.520 24.810 ;
        RECT 258.160 24.490 258.420 24.810 ;
        RECT 258.220 2.400 258.360 24.490 ;
        RECT 258.010 -4.800 258.570 2.400 ;
      LAYER via2 ;
        RECT 21.250 1628.800 21.530 1629.080 ;
      LAYER met3 ;
        RECT 35.000 1631.000 39.000 1631.600 ;
        RECT 21.225 1629.090 21.555 1629.105 ;
        RECT 35.270 1629.090 35.570 1631.000 ;
        RECT 21.225 1628.790 35.570 1629.090 ;
        RECT 21.225 1628.775 21.555 1628.790 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 21.690 24.380 22.010 24.440 ;
        RECT 276.070 24.380 276.390 24.440 ;
        RECT 21.690 24.240 276.390 24.380 ;
        RECT 21.690 24.180 22.010 24.240 ;
        RECT 276.070 24.180 276.390 24.240 ;
      LAYER via ;
        RECT 21.720 24.180 21.980 24.440 ;
        RECT 276.100 24.180 276.360 24.440 ;
      LAYER met2 ;
        RECT 21.710 1732.115 21.990 1732.485 ;
        RECT 21.780 24.470 21.920 1732.115 ;
        RECT 21.720 24.150 21.980 24.470 ;
        RECT 276.100 24.150 276.360 24.470 ;
        RECT 276.160 2.400 276.300 24.150 ;
        RECT 275.950 -4.800 276.510 2.400 ;
      LAYER via2 ;
        RECT 21.710 1732.160 21.990 1732.440 ;
      LAYER met3 ;
        RECT 35.000 1734.360 39.000 1734.960 ;
        RECT 21.685 1732.450 22.015 1732.465 ;
        RECT 35.270 1732.450 35.570 1734.360 ;
        RECT 21.685 1732.150 35.570 1732.450 ;
        RECT 21.685 1732.135 22.015 1732.150 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 48.370 3446.820 48.690 3446.880 ;
        RECT 1459.650 3446.820 1459.970 3446.880 ;
        RECT 48.370 3446.680 1459.970 3446.820 ;
        RECT 48.370 3446.620 48.690 3446.680 ;
        RECT 1459.650 3446.620 1459.970 3446.680 ;
        RECT 48.370 16.220 48.690 16.280 ;
        RECT 294.010 16.220 294.330 16.280 ;
        RECT 48.370 16.080 294.330 16.220 ;
        RECT 48.370 16.020 48.690 16.080 ;
        RECT 294.010 16.020 294.330 16.080 ;
      LAYER via ;
        RECT 48.400 3446.620 48.660 3446.880 ;
        RECT 1459.680 3446.620 1459.940 3446.880 ;
        RECT 48.400 16.020 48.660 16.280 ;
        RECT 294.040 16.020 294.300 16.280 ;
      LAYER met2 ;
        RECT 48.400 3446.590 48.660 3446.910 ;
        RECT 1459.680 3446.590 1459.940 3446.910 ;
        RECT 48.460 16.310 48.600 3446.590 ;
        RECT 1459.740 3435.000 1459.880 3446.590 ;
        RECT 1459.710 3431.000 1459.990 3435.000 ;
        RECT 48.400 15.990 48.660 16.310 ;
        RECT 294.040 15.990 294.300 16.310 ;
        RECT 294.100 2.400 294.240 15.990 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.910 3446.480 48.230 3446.540 ;
        RECT 1564.990 3446.480 1565.310 3446.540 ;
        RECT 47.910 3446.340 1565.310 3446.480 ;
        RECT 47.910 3446.280 48.230 3446.340 ;
        RECT 1564.990 3446.280 1565.310 3446.340 ;
        RECT 47.910 18.260 48.230 18.320 ;
        RECT 311.950 18.260 312.270 18.320 ;
        RECT 47.910 18.120 312.270 18.260 ;
        RECT 47.910 18.060 48.230 18.120 ;
        RECT 311.950 18.060 312.270 18.120 ;
      LAYER via ;
        RECT 47.940 3446.280 48.200 3446.540 ;
        RECT 1565.020 3446.280 1565.280 3446.540 ;
        RECT 47.940 18.060 48.200 18.320 ;
        RECT 311.980 18.060 312.240 18.320 ;
      LAYER met2 ;
        RECT 47.940 3446.250 48.200 3446.570 ;
        RECT 1565.020 3446.250 1565.280 3446.570 ;
        RECT 48.000 18.350 48.140 3446.250 ;
        RECT 1565.080 3435.000 1565.220 3446.250 ;
        RECT 1565.050 3431.000 1565.330 3435.000 ;
        RECT 47.940 18.030 48.200 18.350 ;
        RECT 311.980 18.030 312.240 18.350 ;
        RECT 312.040 2.400 312.180 18.030 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 26.080 330.210 26.140 ;
        RECT 2299.610 26.080 2299.930 26.140 ;
        RECT 329.890 25.940 2299.930 26.080 ;
        RECT 329.890 25.880 330.210 25.940 ;
        RECT 2299.610 25.880 2299.930 25.940 ;
      LAYER via ;
        RECT 329.920 25.880 330.180 26.140 ;
        RECT 2299.640 25.880 2299.900 26.140 ;
      LAYER met2 ;
        RECT 2299.670 35.000 2299.950 39.000 ;
        RECT 2299.700 26.170 2299.840 35.000 ;
        RECT 329.920 25.850 330.180 26.170 ;
        RECT 2299.640 25.850 2299.900 26.170 ;
        RECT 329.980 2.400 330.120 25.850 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 25.740 347.690 25.800 ;
        RECT 2350.210 25.740 2350.530 25.800 ;
        RECT 347.370 25.600 2350.530 25.740 ;
        RECT 347.370 25.540 347.690 25.600 ;
        RECT 2350.210 25.540 2350.530 25.600 ;
      LAYER via ;
        RECT 347.400 25.540 347.660 25.800 ;
        RECT 2350.240 25.540 2350.500 25.800 ;
      LAYER met2 ;
        RECT 2350.270 35.000 2350.550 39.000 ;
        RECT 2350.300 25.830 2350.440 35.000 ;
        RECT 347.400 25.510 347.660 25.830 ;
        RECT 2350.240 25.510 2350.500 25.830 ;
        RECT 347.460 2.400 347.600 25.510 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 24.380 365.630 24.440 ;
        RECT 2401.270 24.380 2401.590 24.440 ;
        RECT 365.310 24.240 2401.590 24.380 ;
        RECT 365.310 24.180 365.630 24.240 ;
        RECT 2401.270 24.180 2401.590 24.240 ;
      LAYER via ;
        RECT 365.340 24.180 365.600 24.440 ;
        RECT 2401.300 24.180 2401.560 24.440 ;
      LAYER met2 ;
        RECT 2401.330 35.000 2401.610 39.000 ;
        RECT 2401.360 24.470 2401.500 35.000 ;
        RECT 365.340 24.150 365.600 24.470 ;
        RECT 2401.300 24.150 2401.560 24.470 ;
        RECT 365.400 2.400 365.540 24.150 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 348.365 16.405 348.535 20.315 ;
      LAYER mcon ;
        RECT 348.365 20.145 348.535 20.315 ;
      LAYER met1 ;
        RECT 45.150 3446.140 45.470 3446.200 ;
        RECT 1670.790 3446.140 1671.110 3446.200 ;
        RECT 45.150 3446.000 1671.110 3446.140 ;
        RECT 45.150 3445.940 45.470 3446.000 ;
        RECT 1670.790 3445.940 1671.110 3446.000 ;
        RECT 45.150 20.300 45.470 20.360 ;
        RECT 348.305 20.300 348.595 20.345 ;
        RECT 45.150 20.160 348.595 20.300 ;
        RECT 45.150 20.100 45.470 20.160 ;
        RECT 348.305 20.115 348.595 20.160 ;
        RECT 348.305 16.560 348.595 16.605 ;
        RECT 383.250 16.560 383.570 16.620 ;
        RECT 348.305 16.420 383.570 16.560 ;
        RECT 348.305 16.375 348.595 16.420 ;
        RECT 383.250 16.360 383.570 16.420 ;
      LAYER via ;
        RECT 45.180 3445.940 45.440 3446.200 ;
        RECT 1670.820 3445.940 1671.080 3446.200 ;
        RECT 45.180 20.100 45.440 20.360 ;
        RECT 383.280 16.360 383.540 16.620 ;
      LAYER met2 ;
        RECT 45.180 3445.910 45.440 3446.230 ;
        RECT 1670.820 3445.910 1671.080 3446.230 ;
        RECT 45.240 20.390 45.380 3445.910 ;
        RECT 1670.880 3435.000 1671.020 3445.910 ;
        RECT 1670.850 3431.000 1671.130 3435.000 ;
        RECT 45.180 20.070 45.440 20.390 ;
        RECT 383.280 16.330 383.540 16.650 ;
        RECT 383.340 2.400 383.480 16.330 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 41.010 3445.800 41.330 3445.860 ;
        RECT 1776.130 3445.800 1776.450 3445.860 ;
        RECT 41.010 3445.660 1776.450 3445.800 ;
        RECT 41.010 3445.600 41.330 3445.660 ;
        RECT 1776.130 3445.600 1776.450 3445.660 ;
        RECT 41.010 19.960 41.330 20.020 ;
        RECT 401.190 19.960 401.510 20.020 ;
        RECT 41.010 19.820 401.510 19.960 ;
        RECT 41.010 19.760 41.330 19.820 ;
        RECT 401.190 19.760 401.510 19.820 ;
      LAYER via ;
        RECT 41.040 3445.600 41.300 3445.860 ;
        RECT 1776.160 3445.600 1776.420 3445.860 ;
        RECT 41.040 19.760 41.300 20.020 ;
        RECT 401.220 19.760 401.480 20.020 ;
      LAYER met2 ;
        RECT 41.040 3445.570 41.300 3445.890 ;
        RECT 1776.160 3445.570 1776.420 3445.890 ;
        RECT 41.100 20.050 41.240 3445.570 ;
        RECT 1776.220 3435.000 1776.360 3445.570 ;
        RECT 1776.190 3431.000 1776.470 3435.000 ;
        RECT 41.040 19.730 41.300 20.050 ;
        RECT 401.220 19.730 401.480 20.050 ;
        RECT 401.280 2.400 401.420 19.730 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2198.010 35.000 2198.290 39.000 ;
        RECT 2198.040 27.725 2198.180 35.000 ;
        RECT 62.190 27.355 62.470 27.725 ;
        RECT 2197.970 27.355 2198.250 27.725 ;
        RECT 62.260 2.400 62.400 27.355 ;
        RECT 62.050 -4.800 62.610 2.400 ;
      LAYER via2 ;
        RECT 62.190 27.400 62.470 27.680 ;
        RECT 2197.970 27.400 2198.250 27.680 ;
      LAYER met3 ;
        RECT 62.165 27.690 62.495 27.705 ;
        RECT 2197.945 27.690 2198.275 27.705 ;
        RECT 62.165 27.390 2198.275 27.690 ;
        RECT 62.165 27.375 62.495 27.390 ;
        RECT 2197.945 27.375 2198.275 27.390 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 24.720 419.450 24.780 ;
        RECT 2452.330 24.720 2452.650 24.780 ;
        RECT 419.130 24.580 2452.650 24.720 ;
        RECT 419.130 24.520 419.450 24.580 ;
        RECT 2452.330 24.520 2452.650 24.580 ;
      LAYER via ;
        RECT 419.160 24.520 419.420 24.780 ;
        RECT 2452.360 24.520 2452.620 24.780 ;
      LAYER met2 ;
        RECT 2452.390 35.000 2452.670 39.000 ;
        RECT 2452.420 24.810 2452.560 35.000 ;
        RECT 419.160 24.490 419.420 24.810 ;
        RECT 2452.360 24.490 2452.620 24.810 ;
        RECT 419.220 2.400 419.360 24.490 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 22.150 30.500 22.470 30.560 ;
        RECT 436.610 30.500 436.930 30.560 ;
        RECT 22.150 30.360 436.930 30.500 ;
        RECT 22.150 30.300 22.470 30.360 ;
        RECT 436.610 30.300 436.930 30.360 ;
      LAYER via ;
        RECT 22.180 30.300 22.440 30.560 ;
        RECT 436.640 30.300 436.900 30.560 ;
      LAYER met2 ;
        RECT 22.170 1836.155 22.450 1836.525 ;
        RECT 22.240 30.590 22.380 1836.155 ;
        RECT 22.180 30.270 22.440 30.590 ;
        RECT 436.640 30.270 436.900 30.590 ;
        RECT 436.700 2.400 436.840 30.270 ;
        RECT 436.490 -4.800 437.050 2.400 ;
      LAYER via2 ;
        RECT 22.170 1836.200 22.450 1836.480 ;
      LAYER met3 ;
        RECT 35.000 1837.040 39.000 1837.640 ;
        RECT 22.145 1836.490 22.475 1836.505 ;
        RECT 35.270 1836.490 35.570 1837.040 ;
        RECT 22.145 1836.190 35.570 1836.490 ;
        RECT 22.145 1836.175 22.475 1836.190 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 22.610 32.880 22.930 32.940 ;
        RECT 454.550 32.880 454.870 32.940 ;
        RECT 22.610 32.740 454.870 32.880 ;
        RECT 22.610 32.680 22.930 32.740 ;
        RECT 454.550 32.680 454.870 32.740 ;
      LAYER via ;
        RECT 22.640 32.680 22.900 32.940 ;
        RECT 454.580 32.680 454.840 32.940 ;
      LAYER met2 ;
        RECT 22.630 1938.835 22.910 1939.205 ;
        RECT 22.700 32.970 22.840 1938.835 ;
        RECT 22.640 32.650 22.900 32.970 ;
        RECT 454.580 32.650 454.840 32.970 ;
        RECT 454.640 2.400 454.780 32.650 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 22.630 1938.880 22.910 1939.160 ;
      LAYER met3 ;
        RECT 35.000 1940.400 39.000 1941.000 ;
        RECT 22.605 1939.170 22.935 1939.185 ;
        RECT 35.270 1939.170 35.570 1940.400 ;
        RECT 22.605 1938.870 35.570 1939.170 ;
        RECT 22.605 1938.855 22.935 1938.870 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 472.490 30.500 472.810 30.560 ;
        RECT 2896.690 30.500 2897.010 30.560 ;
        RECT 472.490 30.360 2897.010 30.500 ;
        RECT 472.490 30.300 472.810 30.360 ;
        RECT 2896.690 30.300 2897.010 30.360 ;
      LAYER via ;
        RECT 472.520 30.300 472.780 30.560 ;
        RECT 2896.720 30.300 2896.980 30.560 ;
      LAYER met2 ;
        RECT 2896.710 1549.195 2896.990 1549.565 ;
        RECT 2896.780 30.590 2896.920 1549.195 ;
        RECT 472.520 30.270 472.780 30.590 ;
        RECT 2896.720 30.270 2896.980 30.590 ;
        RECT 472.580 2.400 472.720 30.270 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 2896.710 1549.240 2896.990 1549.520 ;
      LAYER met3 ;
        RECT 2881.000 1552.120 2885.000 1552.720 ;
        RECT 2884.510 1549.530 2884.810 1552.120 ;
        RECT 2896.685 1549.530 2897.015 1549.545 ;
        RECT 2884.510 1549.230 2897.015 1549.530 ;
        RECT 2896.685 1549.215 2897.015 1549.230 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 490.430 25.400 490.750 25.460 ;
        RECT 2502.930 25.400 2503.250 25.460 ;
        RECT 490.430 25.260 2503.250 25.400 ;
        RECT 490.430 25.200 490.750 25.260 ;
        RECT 2502.930 25.200 2503.250 25.260 ;
      LAYER via ;
        RECT 490.460 25.200 490.720 25.460 ;
        RECT 2502.960 25.200 2503.220 25.460 ;
      LAYER met2 ;
        RECT 2502.990 35.000 2503.270 39.000 ;
        RECT 2503.020 25.490 2503.160 35.000 ;
        RECT 490.460 25.170 490.720 25.490 ;
        RECT 2502.960 25.170 2503.220 25.490 ;
        RECT 490.520 2.400 490.660 25.170 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.070 29.820 23.390 29.880 ;
        RECT 507.910 29.820 508.230 29.880 ;
        RECT 23.070 29.680 508.230 29.820 ;
        RECT 23.070 29.620 23.390 29.680 ;
        RECT 507.910 29.620 508.230 29.680 ;
      LAYER via ;
        RECT 23.100 29.620 23.360 29.880 ;
        RECT 507.940 29.620 508.200 29.880 ;
      LAYER met2 ;
        RECT 23.090 2042.875 23.370 2043.245 ;
        RECT 23.160 29.910 23.300 2042.875 ;
        RECT 23.100 29.590 23.360 29.910 ;
        RECT 507.940 29.590 508.200 29.910 ;
        RECT 508.000 2.400 508.140 29.590 ;
        RECT 507.790 -4.800 508.350 2.400 ;
      LAYER via2 ;
        RECT 23.090 2042.920 23.370 2043.200 ;
      LAYER met3 ;
        RECT 23.065 2043.210 23.395 2043.225 ;
        RECT 35.000 2043.210 39.000 2043.680 ;
        RECT 23.065 2043.080 39.000 2043.210 ;
        RECT 23.065 2042.910 35.570 2043.080 ;
        RECT 23.065 2042.895 23.395 2042.910 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.530 30.160 23.850 30.220 ;
        RECT 525.850 30.160 526.170 30.220 ;
        RECT 23.530 30.020 526.170 30.160 ;
        RECT 23.530 29.960 23.850 30.020 ;
        RECT 525.850 29.960 526.170 30.020 ;
      LAYER via ;
        RECT 23.560 29.960 23.820 30.220 ;
        RECT 525.880 29.960 526.140 30.220 ;
      LAYER met2 ;
        RECT 23.550 2146.235 23.830 2146.605 ;
        RECT 23.620 30.250 23.760 2146.235 ;
        RECT 23.560 29.930 23.820 30.250 ;
        RECT 525.880 29.930 526.140 30.250 ;
        RECT 525.940 2.400 526.080 29.930 ;
        RECT 525.730 -4.800 526.290 2.400 ;
      LAYER via2 ;
        RECT 23.550 2146.280 23.830 2146.560 ;
      LAYER met3 ;
        RECT 23.525 2146.570 23.855 2146.585 ;
        RECT 35.000 2146.570 39.000 2147.040 ;
        RECT 23.525 2146.440 39.000 2146.570 ;
        RECT 23.525 2146.270 35.570 2146.440 ;
        RECT 23.525 2146.255 23.855 2146.270 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 543.790 30.160 544.110 30.220 ;
        RECT 2896.230 30.160 2896.550 30.220 ;
        RECT 543.790 30.020 2896.550 30.160 ;
        RECT 543.790 29.960 544.110 30.020 ;
        RECT 2896.230 29.960 2896.550 30.020 ;
      LAYER via ;
        RECT 543.820 29.960 544.080 30.220 ;
        RECT 2896.260 29.960 2896.520 30.220 ;
      LAYER met2 ;
        RECT 2896.250 1670.915 2896.530 1671.285 ;
        RECT 2896.320 30.250 2896.460 1670.915 ;
        RECT 543.820 29.930 544.080 30.250 ;
        RECT 2896.260 29.930 2896.520 30.250 ;
        RECT 543.880 2.400 544.020 29.930 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 2896.250 1670.960 2896.530 1671.240 ;
      LAYER met3 ;
        RECT 2881.000 1673.840 2885.000 1674.440 ;
        RECT 2884.510 1671.250 2884.810 1673.840 ;
        RECT 2896.225 1671.250 2896.555 1671.265 ;
        RECT 2884.510 1670.950 2896.555 1671.250 ;
        RECT 2896.225 1670.935 2896.555 1670.950 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 29.820 562.050 29.880 ;
        RECT 2895.770 29.820 2896.090 29.880 ;
        RECT 561.730 29.680 2896.090 29.820 ;
        RECT 561.730 29.620 562.050 29.680 ;
        RECT 2895.770 29.620 2896.090 29.680 ;
      LAYER via ;
        RECT 561.760 29.620 562.020 29.880 ;
        RECT 2895.800 29.620 2896.060 29.880 ;
      LAYER met2 ;
        RECT 2895.790 1793.995 2896.070 1794.365 ;
        RECT 2895.860 29.910 2896.000 1793.995 ;
        RECT 561.760 29.590 562.020 29.910 ;
        RECT 2895.800 29.590 2896.060 29.910 ;
        RECT 561.820 2.400 561.960 29.590 ;
        RECT 561.610 -4.800 562.170 2.400 ;
      LAYER via2 ;
        RECT 2895.790 1794.040 2896.070 1794.320 ;
      LAYER met3 ;
        RECT 2881.000 1795.560 2885.000 1796.160 ;
        RECT 2884.510 1794.330 2884.810 1795.560 ;
        RECT 2895.765 1794.330 2896.095 1794.345 ;
        RECT 2884.510 1794.030 2896.095 1794.330 ;
        RECT 2895.765 1794.015 2896.095 1794.030 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.990 29.480 24.310 29.540 ;
        RECT 579.670 29.480 579.990 29.540 ;
        RECT 23.990 29.340 579.990 29.480 ;
        RECT 23.990 29.280 24.310 29.340 ;
        RECT 579.670 29.280 579.990 29.340 ;
      LAYER via ;
        RECT 24.020 29.280 24.280 29.540 ;
        RECT 579.700 29.280 579.960 29.540 ;
      LAYER met2 ;
        RECT 24.010 2249.595 24.290 2249.965 ;
        RECT 24.080 29.570 24.220 2249.595 ;
        RECT 24.020 29.250 24.280 29.570 ;
        RECT 579.700 29.250 579.960 29.570 ;
        RECT 579.760 2.400 579.900 29.250 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 24.010 2249.640 24.290 2249.920 ;
      LAYER met3 ;
        RECT 23.985 2249.930 24.315 2249.945 ;
        RECT 23.985 2249.720 35.570 2249.930 ;
        RECT 23.985 2249.630 39.000 2249.720 ;
        RECT 23.985 2249.615 24.315 2249.630 ;
        RECT 35.000 2249.120 39.000 2249.630 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 40.550 3447.500 40.870 3447.560 ;
        RECT 1248.510 3447.500 1248.830 3447.560 ;
        RECT 40.550 3447.360 1248.830 3447.500 ;
        RECT 40.550 3447.300 40.870 3447.360 ;
        RECT 1248.510 3447.300 1248.830 3447.360 ;
        RECT 40.550 14.180 40.870 14.240 ;
        RECT 86.090 14.180 86.410 14.240 ;
        RECT 40.550 14.040 86.410 14.180 ;
        RECT 40.550 13.980 40.870 14.040 ;
        RECT 86.090 13.980 86.410 14.040 ;
      LAYER via ;
        RECT 40.580 3447.300 40.840 3447.560 ;
        RECT 1248.540 3447.300 1248.800 3447.560 ;
        RECT 40.580 13.980 40.840 14.240 ;
        RECT 86.120 13.980 86.380 14.240 ;
      LAYER met2 ;
        RECT 40.580 3447.270 40.840 3447.590 ;
        RECT 1248.540 3447.270 1248.800 3447.590 ;
        RECT 40.640 14.270 40.780 3447.270 ;
        RECT 1248.600 3435.000 1248.740 3447.270 ;
        RECT 1248.570 3431.000 1248.850 3435.000 ;
        RECT 40.580 13.950 40.840 14.270 ;
        RECT 86.120 13.950 86.380 14.270 ;
        RECT 86.180 2.400 86.320 13.950 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 597.150 29.480 597.470 29.540 ;
        RECT 2895.310 29.480 2895.630 29.540 ;
        RECT 597.150 29.340 2895.630 29.480 ;
        RECT 597.150 29.280 597.470 29.340 ;
        RECT 2895.310 29.280 2895.630 29.340 ;
      LAYER via ;
        RECT 597.180 29.280 597.440 29.540 ;
        RECT 2895.340 29.280 2895.600 29.540 ;
      LAYER met2 ;
        RECT 2895.330 1913.675 2895.610 1914.045 ;
        RECT 2895.400 29.570 2895.540 1913.675 ;
        RECT 597.180 29.250 597.440 29.570 ;
        RECT 2895.340 29.250 2895.600 29.570 ;
        RECT 597.240 2.400 597.380 29.250 ;
        RECT 597.030 -4.800 597.590 2.400 ;
      LAYER via2 ;
        RECT 2895.330 1913.720 2895.610 1914.000 ;
      LAYER met3 ;
        RECT 2881.000 1916.600 2885.000 1917.200 ;
        RECT 2884.510 1914.010 2884.810 1916.600 ;
        RECT 2895.305 1914.010 2895.635 1914.025 ;
        RECT 2884.510 1913.710 2895.635 1914.010 ;
        RECT 2895.305 1913.695 2895.635 1913.710 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.450 29.140 24.770 29.200 ;
        RECT 615.090 29.140 615.410 29.200 ;
        RECT 24.450 29.000 615.410 29.140 ;
        RECT 24.450 28.940 24.770 29.000 ;
        RECT 615.090 28.940 615.410 29.000 ;
      LAYER via ;
        RECT 24.480 28.940 24.740 29.200 ;
        RECT 615.120 28.940 615.380 29.200 ;
      LAYER met2 ;
        RECT 24.470 2349.555 24.750 2349.925 ;
        RECT 24.540 29.230 24.680 2349.555 ;
        RECT 24.480 28.910 24.740 29.230 ;
        RECT 615.120 28.910 615.380 29.230 ;
        RECT 615.180 2.400 615.320 28.910 ;
        RECT 614.970 -4.800 615.530 2.400 ;
      LAYER via2 ;
        RECT 24.470 2349.600 24.750 2349.880 ;
      LAYER met3 ;
        RECT 35.000 2352.480 39.000 2353.080 ;
        RECT 24.445 2349.890 24.775 2349.905 ;
        RECT 35.270 2349.890 35.570 2352.480 ;
        RECT 24.445 2349.590 35.570 2349.890 ;
        RECT 24.445 2349.575 24.775 2349.590 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 46.070 3447.160 46.390 3447.220 ;
        RECT 1353.850 3447.160 1354.170 3447.220 ;
        RECT 46.070 3447.020 1354.170 3447.160 ;
        RECT 46.070 3446.960 46.390 3447.020 ;
        RECT 1353.850 3446.960 1354.170 3447.020 ;
        RECT 46.070 14.520 46.390 14.580 ;
        RECT 109.550 14.520 109.870 14.580 ;
        RECT 46.070 14.380 109.870 14.520 ;
        RECT 46.070 14.320 46.390 14.380 ;
        RECT 109.550 14.320 109.870 14.380 ;
      LAYER via ;
        RECT 46.100 3446.960 46.360 3447.220 ;
        RECT 1353.880 3446.960 1354.140 3447.220 ;
        RECT 46.100 14.320 46.360 14.580 ;
        RECT 109.580 14.320 109.840 14.580 ;
      LAYER met2 ;
        RECT 46.100 3446.930 46.360 3447.250 ;
        RECT 1353.880 3446.930 1354.140 3447.250 ;
        RECT 46.160 14.610 46.300 3446.930 ;
        RECT 1353.940 3435.000 1354.080 3446.930 ;
        RECT 1353.910 3431.000 1354.190 3435.000 ;
        RECT 46.100 14.290 46.360 14.610 ;
        RECT 109.580 14.290 109.840 14.610 ;
        RECT 109.640 2.400 109.780 14.290 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.730 17.240 33.050 17.300 ;
        RECT 133.470 17.240 133.790 17.300 ;
        RECT 32.730 17.100 133.790 17.240 ;
        RECT 32.730 17.040 33.050 17.100 ;
        RECT 133.470 17.040 133.790 17.100 ;
      LAYER via ;
        RECT 32.760 17.040 33.020 17.300 ;
        RECT 133.500 17.040 133.760 17.300 ;
      LAYER met2 ;
        RECT 32.750 1218.035 33.030 1218.405 ;
        RECT 32.820 17.330 32.960 1218.035 ;
        RECT 32.760 17.010 33.020 17.330 ;
        RECT 133.500 17.010 133.760 17.330 ;
        RECT 133.560 2.400 133.700 17.010 ;
        RECT 133.350 -4.800 133.910 2.400 ;
      LAYER via2 ;
        RECT 32.750 1218.080 33.030 1218.360 ;
      LAYER met3 ;
        RECT 35.000 1218.920 39.000 1219.520 ;
        RECT 32.725 1218.370 33.055 1218.385 ;
        RECT 35.270 1218.370 35.570 1218.920 ;
        RECT 32.725 1218.070 35.570 1218.370 ;
        RECT 32.725 1218.055 33.055 1218.070 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 30.840 151.730 30.900 ;
        RECT 2897.610 30.840 2897.930 30.900 ;
        RECT 151.410 30.700 2897.930 30.840 ;
        RECT 151.410 30.640 151.730 30.700 ;
        RECT 2897.610 30.640 2897.930 30.700 ;
      LAYER via ;
        RECT 151.440 30.640 151.700 30.900 ;
        RECT 2897.640 30.640 2897.900 30.900 ;
      LAYER met2 ;
        RECT 2897.630 1306.435 2897.910 1306.805 ;
        RECT 2897.700 30.930 2897.840 1306.435 ;
        RECT 151.440 30.610 151.700 30.930 ;
        RECT 2897.640 30.610 2897.900 30.930 ;
        RECT 151.500 2.400 151.640 30.610 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 2897.630 1306.480 2897.910 1306.760 ;
      LAYER met3 ;
        RECT 2881.000 1309.360 2885.000 1309.960 ;
        RECT 2884.510 1306.770 2884.810 1309.360 ;
        RECT 2897.605 1306.770 2897.935 1306.785 ;
        RECT 2884.510 1306.470 2897.935 1306.770 ;
        RECT 2897.605 1306.455 2897.935 1306.470 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 169.350 31.180 169.670 31.240 ;
        RECT 2897.150 31.180 2897.470 31.240 ;
        RECT 169.350 31.040 2897.470 31.180 ;
        RECT 169.350 30.980 169.670 31.040 ;
        RECT 2897.150 30.980 2897.470 31.040 ;
      LAYER via ;
        RECT 169.380 30.980 169.640 31.240 ;
        RECT 2897.180 30.980 2897.440 31.240 ;
      LAYER met2 ;
        RECT 2897.170 1428.155 2897.450 1428.525 ;
        RECT 2897.240 31.270 2897.380 1428.155 ;
        RECT 169.380 30.950 169.640 31.270 ;
        RECT 2897.180 30.950 2897.440 31.270 ;
        RECT 169.440 2.400 169.580 30.950 ;
        RECT 169.230 -4.800 169.790 2.400 ;
      LAYER via2 ;
        RECT 2897.170 1428.200 2897.450 1428.480 ;
      LAYER met3 ;
        RECT 2881.000 1431.080 2885.000 1431.680 ;
        RECT 2884.510 1428.490 2884.810 1431.080 ;
        RECT 2897.145 1428.490 2897.475 1428.505 ;
        RECT 2884.510 1428.190 2897.475 1428.490 ;
        RECT 2897.145 1428.175 2897.475 1428.190 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 35.490 14.860 35.810 14.920 ;
        RECT 186.830 14.860 187.150 14.920 ;
        RECT 35.490 14.720 187.150 14.860 ;
        RECT 35.490 14.660 35.810 14.720 ;
        RECT 186.830 14.660 187.150 14.720 ;
      LAYER via ;
        RECT 35.520 14.660 35.780 14.920 ;
        RECT 186.860 14.660 187.120 14.920 ;
      LAYER met2 ;
        RECT 35.510 1319.355 35.790 1319.725 ;
        RECT 35.580 14.950 35.720 1319.355 ;
        RECT 35.520 14.630 35.780 14.950 ;
        RECT 186.860 14.630 187.120 14.950 ;
        RECT 186.920 2.400 187.060 14.630 ;
        RECT 186.710 -4.800 187.270 2.400 ;
      LAYER via2 ;
        RECT 35.510 1319.400 35.790 1319.680 ;
      LAYER met3 ;
        RECT 35.000 1322.280 39.000 1322.880 ;
        RECT 35.270 1319.705 35.570 1322.280 ;
        RECT 35.270 1319.390 35.815 1319.705 ;
        RECT 35.485 1319.375 35.815 1319.390 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 33.190 15.200 33.510 15.260 ;
        RECT 204.770 15.200 205.090 15.260 ;
        RECT 33.190 15.060 205.090 15.200 ;
        RECT 33.190 15.000 33.510 15.060 ;
        RECT 204.770 15.000 205.090 15.060 ;
      LAYER via ;
        RECT 33.220 15.000 33.480 15.260 ;
        RECT 204.800 15.000 205.060 15.260 ;
      LAYER met2 ;
        RECT 33.210 1424.075 33.490 1424.445 ;
        RECT 33.280 15.290 33.420 1424.075 ;
        RECT 33.220 14.970 33.480 15.290 ;
        RECT 204.800 14.970 205.060 15.290 ;
        RECT 204.860 2.400 205.000 14.970 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 33.210 1424.120 33.490 1424.400 ;
      LAYER met3 ;
        RECT 35.000 1424.960 39.000 1425.560 ;
        RECT 33.185 1424.410 33.515 1424.425 ;
        RECT 35.270 1424.410 35.570 1424.960 ;
        RECT 33.185 1424.110 35.570 1424.410 ;
        RECT 33.185 1424.095 33.515 1424.110 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 35.030 15.540 35.350 15.600 ;
        RECT 222.710 15.540 223.030 15.600 ;
        RECT 35.030 15.400 223.030 15.540 ;
        RECT 35.030 15.340 35.350 15.400 ;
        RECT 222.710 15.340 223.030 15.400 ;
      LAYER via ;
        RECT 35.060 15.340 35.320 15.600 ;
        RECT 222.740 15.340 223.000 15.600 ;
      LAYER met2 ;
        RECT 35.050 1525.395 35.330 1525.765 ;
        RECT 35.120 15.630 35.260 1525.395 ;
        RECT 35.060 15.310 35.320 15.630 ;
        RECT 222.740 15.310 223.000 15.630 ;
        RECT 222.800 2.400 222.940 15.310 ;
        RECT 222.590 -4.800 223.150 2.400 ;
      LAYER via2 ;
        RECT 35.050 1525.440 35.330 1525.720 ;
      LAYER met3 ;
        RECT 35.000 1528.320 39.000 1528.920 ;
        RECT 35.270 1525.745 35.570 1528.320 ;
        RECT 35.025 1525.430 35.570 1525.745 ;
        RECT 35.025 1525.415 35.355 1525.430 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 3445.120 20.630 3445.180 ;
        RECT 1881.930 3445.120 1882.250 3445.180 ;
        RECT 20.310 3444.980 1882.250 3445.120 ;
        RECT 20.310 3444.920 20.630 3444.980 ;
        RECT 1881.930 3444.920 1882.250 3444.980 ;
      LAYER via ;
        RECT 20.340 3444.920 20.600 3445.180 ;
        RECT 1881.960 3444.920 1882.220 3445.180 ;
      LAYER met2 ;
        RECT 20.340 3444.890 20.600 3445.210 ;
        RECT 1881.960 3444.890 1882.220 3445.210 ;
        RECT 20.400 2.400 20.540 3444.890 ;
        RECT 1882.020 3435.000 1882.160 3444.890 ;
        RECT 1881.990 3431.000 1882.270 3435.000 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.910 20.300 25.230 20.360 ;
        RECT 44.230 20.300 44.550 20.360 ;
        RECT 24.910 20.160 44.550 20.300 ;
        RECT 24.910 20.100 25.230 20.160 ;
        RECT 44.230 20.100 44.550 20.160 ;
      LAYER via ;
        RECT 24.940 20.100 25.200 20.360 ;
        RECT 44.260 20.100 44.520 20.360 ;
      LAYER met2 ;
        RECT 24.930 2452.235 25.210 2452.605 ;
        RECT 25.000 20.390 25.140 2452.235 ;
        RECT 24.940 20.070 25.200 20.390 ;
        RECT 44.260 20.070 44.520 20.390 ;
        RECT 44.320 2.400 44.460 20.070 ;
        RECT 44.110 -4.800 44.670 2.400 ;
      LAYER via2 ;
        RECT 24.930 2452.280 25.210 2452.560 ;
      LAYER met3 ;
        RECT 35.000 2455.160 39.000 2455.760 ;
        RECT 24.905 2452.570 25.235 2452.585 ;
        RECT 35.270 2452.570 35.570 2455.160 ;
        RECT 24.905 2452.270 35.570 2452.570 ;
        RECT 24.905 2452.255 25.235 2452.270 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 33.650 16.900 33.970 16.960 ;
        RECT 246.630 16.900 246.950 16.960 ;
        RECT 33.650 16.760 246.950 16.900 ;
        RECT 33.650 16.700 33.970 16.760 ;
        RECT 246.630 16.700 246.950 16.760 ;
      LAYER via ;
        RECT 33.680 16.700 33.940 16.960 ;
        RECT 246.660 16.700 246.920 16.960 ;
      LAYER met2 ;
        RECT 33.670 2660.315 33.950 2660.685 ;
        RECT 33.740 16.990 33.880 2660.315 ;
        RECT 33.680 16.670 33.940 16.990 ;
        RECT 246.660 16.670 246.920 16.990 ;
        RECT 246.720 2.400 246.860 16.670 ;
        RECT 246.510 -4.800 247.070 2.400 ;
      LAYER via2 ;
        RECT 33.670 2660.360 33.950 2660.640 ;
      LAYER met3 ;
        RECT 35.000 2661.670 39.000 2661.800 ;
        RECT 33.430 2661.370 39.000 2661.670 ;
        RECT 33.430 2660.665 33.730 2661.370 ;
        RECT 35.000 2661.200 39.000 2661.370 ;
        RECT 33.430 2660.350 33.975 2660.665 ;
        RECT 33.645 2660.335 33.975 2660.350 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 264.110 31.520 264.430 31.580 ;
        RECT 2893.470 31.520 2893.790 31.580 ;
        RECT 264.110 31.380 2893.790 31.520 ;
        RECT 264.110 31.320 264.430 31.380 ;
        RECT 2893.470 31.320 2893.790 31.380 ;
      LAYER via ;
        RECT 264.140 31.320 264.400 31.580 ;
        RECT 2893.500 31.320 2893.760 31.580 ;
      LAYER met2 ;
        RECT 2893.490 2401.915 2893.770 2402.285 ;
        RECT 2893.560 31.610 2893.700 2401.915 ;
        RECT 264.140 31.290 264.400 31.610 ;
        RECT 2893.500 31.290 2893.760 31.610 ;
        RECT 264.200 2.400 264.340 31.290 ;
        RECT 263.990 -4.800 264.550 2.400 ;
      LAYER via2 ;
        RECT 2893.490 2401.960 2893.770 2402.240 ;
      LAYER met3 ;
        RECT 2881.000 2402.250 2885.000 2402.720 ;
        RECT 2893.465 2402.250 2893.795 2402.265 ;
        RECT 2881.000 2402.120 2893.795 2402.250 ;
        RECT 2884.510 2401.950 2893.795 2402.120 ;
        RECT 2893.465 2401.935 2893.795 2401.950 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 31.860 282.370 31.920 ;
        RECT 2893.010 31.860 2893.330 31.920 ;
        RECT 282.050 31.720 2893.330 31.860 ;
        RECT 282.050 31.660 282.370 31.720 ;
        RECT 2893.010 31.660 2893.330 31.720 ;
      LAYER via ;
        RECT 282.080 31.660 282.340 31.920 ;
        RECT 2893.040 31.660 2893.300 31.920 ;
      LAYER met2 ;
        RECT 2893.030 2520.915 2893.310 2521.285 ;
        RECT 2893.100 31.950 2893.240 2520.915 ;
        RECT 282.080 31.630 282.340 31.950 ;
        RECT 2893.040 31.630 2893.300 31.950 ;
        RECT 282.140 2.400 282.280 31.630 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 2893.030 2520.960 2893.310 2521.240 ;
      LAYER met3 ;
        RECT 2881.000 2523.840 2885.000 2524.440 ;
        RECT 2884.510 2521.250 2884.810 2523.840 ;
        RECT 2893.005 2521.250 2893.335 2521.265 ;
        RECT 2884.510 2520.950 2893.335 2521.250 ;
        RECT 2893.005 2520.935 2893.335 2520.950 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 45.610 3444.100 45.930 3444.160 ;
        RECT 2198.410 3444.100 2198.730 3444.160 ;
        RECT 45.610 3443.960 2198.730 3444.100 ;
        RECT 45.610 3443.900 45.930 3443.960 ;
        RECT 2198.410 3443.900 2198.730 3443.960 ;
        RECT 45.610 16.560 45.930 16.620 ;
        RECT 299.990 16.560 300.310 16.620 ;
        RECT 45.610 16.420 300.310 16.560 ;
        RECT 45.610 16.360 45.930 16.420 ;
        RECT 299.990 16.360 300.310 16.420 ;
      LAYER via ;
        RECT 45.640 3443.900 45.900 3444.160 ;
        RECT 2198.440 3443.900 2198.700 3444.160 ;
        RECT 45.640 16.360 45.900 16.620 ;
        RECT 300.020 16.360 300.280 16.620 ;
      LAYER met2 ;
        RECT 45.640 3443.870 45.900 3444.190 ;
        RECT 2198.440 3443.870 2198.700 3444.190 ;
        RECT 45.700 16.650 45.840 3443.870 ;
        RECT 2198.500 3435.000 2198.640 3443.870 ;
        RECT 2198.470 3431.000 2198.750 3435.000 ;
        RECT 45.640 16.330 45.900 16.650 ;
        RECT 300.020 16.330 300.280 16.650 ;
        RECT 300.080 2.400 300.220 16.330 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.930 18.260 318.250 18.320 ;
        RECT 2706.710 18.260 2707.030 18.320 ;
        RECT 317.930 18.120 2707.030 18.260 ;
        RECT 317.930 18.060 318.250 18.120 ;
        RECT 2706.710 18.060 2707.030 18.120 ;
      LAYER via ;
        RECT 317.960 18.060 318.220 18.320 ;
        RECT 2706.740 18.060 2707.000 18.320 ;
      LAYER met2 ;
        RECT 2706.770 35.000 2707.050 39.000 ;
        RECT 2706.800 18.350 2706.940 35.000 ;
        RECT 317.960 18.030 318.220 18.350 ;
        RECT 2706.740 18.030 2707.000 18.350 ;
        RECT 318.020 2.400 318.160 18.030 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 46.990 3443.760 47.310 3443.820 ;
        RECT 2304.210 3443.760 2304.530 3443.820 ;
        RECT 46.990 3443.620 2304.530 3443.760 ;
        RECT 46.990 3443.560 47.310 3443.620 ;
        RECT 2304.210 3443.560 2304.530 3443.620 ;
      LAYER via ;
        RECT 47.020 3443.560 47.280 3443.820 ;
        RECT 2304.240 3443.560 2304.500 3443.820 ;
      LAYER met2 ;
        RECT 47.020 3443.530 47.280 3443.850 ;
        RECT 2304.240 3443.530 2304.500 3443.850 ;
        RECT 47.080 20.245 47.220 3443.530 ;
        RECT 2304.300 3435.000 2304.440 3443.530 ;
        RECT 2304.270 3431.000 2304.550 3435.000 ;
        RECT 47.010 19.875 47.290 20.245 ;
        RECT 335.890 19.875 336.170 20.245 ;
        RECT 335.960 2.400 336.100 19.875 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 47.010 19.920 47.290 20.200 ;
        RECT 335.890 19.920 336.170 20.200 ;
      LAYER met3 ;
        RECT 46.985 20.210 47.315 20.225 ;
        RECT 335.865 20.210 336.195 20.225 ;
        RECT 46.985 19.910 336.195 20.210 ;
        RECT 46.985 19.895 47.315 19.910 ;
        RECT 335.865 19.895 336.195 19.910 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 34.570 20.640 34.890 20.700 ;
        RECT 353.350 20.640 353.670 20.700 ;
        RECT 34.570 20.500 353.670 20.640 ;
        RECT 34.570 20.440 34.890 20.500 ;
        RECT 353.350 20.440 353.670 20.500 ;
      LAYER via ;
        RECT 34.600 20.440 34.860 20.700 ;
        RECT 353.380 20.440 353.640 20.700 ;
      LAYER met2 ;
        RECT 34.590 2761.635 34.870 2762.005 ;
        RECT 34.660 20.730 34.800 2761.635 ;
        RECT 34.600 20.410 34.860 20.730 ;
        RECT 353.380 20.410 353.640 20.730 ;
        RECT 353.440 2.400 353.580 20.410 ;
        RECT 353.230 -4.800 353.790 2.400 ;
      LAYER via2 ;
        RECT 34.590 2761.680 34.870 2761.960 ;
      LAYER met3 ;
        RECT 35.000 2764.560 39.000 2765.160 ;
        RECT 34.565 2761.970 34.895 2761.985 ;
        RECT 35.270 2761.970 35.570 2764.560 ;
        RECT 34.565 2761.670 35.570 2761.970 ;
        RECT 34.565 2761.655 34.895 2761.670 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.450 3443.420 47.770 3443.480 ;
        RECT 2409.550 3443.420 2409.870 3443.480 ;
        RECT 47.450 3443.280 2409.870 3443.420 ;
        RECT 47.450 3443.220 47.770 3443.280 ;
        RECT 2409.550 3443.220 2409.870 3443.280 ;
      LAYER via ;
        RECT 47.480 3443.220 47.740 3443.480 ;
        RECT 2409.580 3443.220 2409.840 3443.480 ;
      LAYER met2 ;
        RECT 47.480 3443.190 47.740 3443.510 ;
        RECT 2409.580 3443.190 2409.840 3443.510 ;
        RECT 47.540 19.565 47.680 3443.190 ;
        RECT 2409.640 3435.000 2409.780 3443.190 ;
        RECT 2409.610 3431.000 2409.890 3435.000 ;
        RECT 47.470 19.195 47.750 19.565 ;
        RECT 371.310 19.195 371.590 19.565 ;
        RECT 371.380 2.400 371.520 19.195 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 47.470 19.240 47.750 19.520 ;
        RECT 371.310 19.240 371.590 19.520 ;
      LAYER met3 ;
        RECT 47.445 19.530 47.775 19.545 ;
        RECT 371.285 19.530 371.615 19.545 ;
        RECT 47.445 19.230 371.615 19.530 ;
        RECT 47.445 19.215 47.775 19.230 ;
        RECT 371.285 19.215 371.615 19.230 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2515.370 3445.035 2515.650 3445.405 ;
        RECT 2515.440 3435.000 2515.580 3445.035 ;
        RECT 2515.410 3431.000 2515.690 3435.000 ;
        RECT 389.250 19.195 389.530 19.565 ;
        RECT 389.320 2.400 389.460 19.195 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 2515.370 3445.080 2515.650 3445.360 ;
        RECT 389.250 19.240 389.530 19.520 ;
      LAYER met3 ;
        RECT 2515.345 3445.370 2515.675 3445.385 ;
        RECT 2849.510 3445.370 2849.890 3445.380 ;
        RECT 2515.345 3445.070 2849.890 3445.370 ;
        RECT 2515.345 3445.055 2515.675 3445.070 ;
        RECT 2849.510 3445.060 2849.890 3445.070 ;
        RECT 389.225 19.530 389.555 19.545 ;
        RECT 2849.510 19.530 2849.890 19.540 ;
        RECT 389.225 19.230 2849.890 19.530 ;
        RECT 389.225 19.215 389.555 19.230 ;
        RECT 2849.510 19.220 2849.890 19.230 ;
      LAYER via3 ;
        RECT 2849.540 3445.060 2849.860 3445.380 ;
        RECT 2849.540 19.220 2849.860 19.540 ;
      LAYER met4 ;
        RECT 2849.535 3445.055 2849.865 3445.385 ;
        RECT 2849.550 19.545 2849.850 3445.055 ;
        RECT 2849.535 19.215 2849.865 19.545 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 407.170 32.200 407.490 32.260 ;
        RECT 2892.550 32.200 2892.870 32.260 ;
        RECT 407.170 32.060 2892.870 32.200 ;
        RECT 407.170 32.000 407.490 32.060 ;
        RECT 2892.550 32.000 2892.870 32.060 ;
      LAYER via ;
        RECT 407.200 32.000 407.460 32.260 ;
        RECT 2892.580 32.000 2892.840 32.260 ;
      LAYER met2 ;
        RECT 2892.570 2643.995 2892.850 2644.365 ;
        RECT 2892.640 32.290 2892.780 2643.995 ;
        RECT 407.200 31.970 407.460 32.290 ;
        RECT 2892.580 31.970 2892.840 32.290 ;
        RECT 407.260 2.400 407.400 31.970 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 2892.570 2644.040 2892.850 2644.320 ;
      LAYER met3 ;
        RECT 2881.000 2645.560 2885.000 2646.160 ;
        RECT 2884.510 2644.330 2884.810 2645.560 ;
        RECT 2892.545 2644.330 2892.875 2644.345 ;
        RECT 2884.510 2644.030 2892.875 2644.330 ;
        RECT 2892.545 2644.015 2892.875 2644.030 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.150 17.920 68.470 17.980 ;
        RECT 2553.990 17.920 2554.310 17.980 ;
        RECT 68.150 17.780 2554.310 17.920 ;
        RECT 68.150 17.720 68.470 17.780 ;
        RECT 2553.990 17.720 2554.310 17.780 ;
      LAYER via ;
        RECT 68.180 17.720 68.440 17.980 ;
        RECT 2554.020 17.720 2554.280 17.980 ;
      LAYER met2 ;
        RECT 2554.050 35.000 2554.330 39.000 ;
        RECT 2554.080 18.010 2554.220 35.000 ;
        RECT 68.180 17.690 68.440 18.010 ;
        RECT 2554.020 17.690 2554.280 18.010 ;
        RECT 68.240 2.400 68.380 17.690 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 424.650 32.540 424.970 32.600 ;
        RECT 2892.090 32.540 2892.410 32.600 ;
        RECT 424.650 32.400 2892.410 32.540 ;
        RECT 424.650 32.340 424.970 32.400 ;
        RECT 2892.090 32.340 2892.410 32.400 ;
      LAYER via ;
        RECT 424.680 32.340 424.940 32.600 ;
        RECT 2892.120 32.340 2892.380 32.600 ;
      LAYER met2 ;
        RECT 2892.110 2767.075 2892.390 2767.445 ;
        RECT 2892.180 32.630 2892.320 2767.075 ;
        RECT 424.680 32.310 424.940 32.630 ;
        RECT 2892.120 32.310 2892.380 32.630 ;
        RECT 424.740 2.400 424.880 32.310 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 2892.110 2767.120 2892.390 2767.400 ;
      LAYER met3 ;
        RECT 2892.085 2767.410 2892.415 2767.425 ;
        RECT 2884.510 2767.200 2892.415 2767.410 ;
        RECT 2881.000 2767.110 2892.415 2767.200 ;
        RECT 2881.000 2766.600 2885.000 2767.110 ;
        RECT 2892.085 2767.095 2892.415 2767.110 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 34.110 19.620 34.430 19.680 ;
        RECT 442.590 19.620 442.910 19.680 ;
        RECT 34.110 19.480 442.910 19.620 ;
        RECT 34.110 19.420 34.430 19.480 ;
        RECT 442.590 19.420 442.910 19.480 ;
      LAYER via ;
        RECT 34.140 19.420 34.400 19.680 ;
        RECT 442.620 19.420 442.880 19.680 ;
      LAYER met2 ;
        RECT 34.130 2866.355 34.410 2866.725 ;
        RECT 34.200 19.710 34.340 2866.355 ;
        RECT 34.140 19.390 34.400 19.710 ;
        RECT 442.620 19.390 442.880 19.710 ;
        RECT 442.680 2.400 442.820 19.390 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 34.130 2866.400 34.410 2866.680 ;
      LAYER met3 ;
        RECT 35.000 2867.240 39.000 2867.840 ;
        RECT 34.105 2866.690 34.435 2866.705 ;
        RECT 35.270 2866.690 35.570 2867.240 ;
        RECT 34.105 2866.390 35.570 2866.690 ;
        RECT 34.105 2866.375 34.435 2866.390 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 460.530 32.880 460.850 32.940 ;
        RECT 2891.630 32.880 2891.950 32.940 ;
        RECT 460.530 32.740 2891.950 32.880 ;
        RECT 460.530 32.680 460.850 32.740 ;
        RECT 2891.630 32.680 2891.950 32.740 ;
      LAYER via ;
        RECT 460.560 32.680 460.820 32.940 ;
        RECT 2891.660 32.680 2891.920 32.940 ;
      LAYER met2 ;
        RECT 2891.650 2886.075 2891.930 2886.445 ;
        RECT 2891.720 32.970 2891.860 2886.075 ;
        RECT 460.560 32.650 460.820 32.970 ;
        RECT 2891.660 32.650 2891.920 32.970 ;
        RECT 460.620 2.400 460.760 32.650 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 2891.650 2886.120 2891.930 2886.400 ;
      LAYER met3 ;
        RECT 2881.000 2888.320 2885.000 2888.920 ;
        RECT 2884.510 2886.410 2884.810 2888.320 ;
        RECT 2891.625 2886.410 2891.955 2886.425 ;
        RECT 2884.510 2886.110 2891.955 2886.410 ;
        RECT 2891.625 2886.095 2891.955 2886.110 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2891.190 3008.475 2891.470 3008.845 ;
        RECT 2891.260 20.245 2891.400 3008.475 ;
        RECT 478.490 19.875 478.770 20.245 ;
        RECT 2891.190 19.875 2891.470 20.245 ;
        RECT 478.560 2.400 478.700 19.875 ;
        RECT 478.350 -4.800 478.910 2.400 ;
      LAYER via2 ;
        RECT 2891.190 3008.520 2891.470 3008.800 ;
        RECT 478.490 19.920 478.770 20.200 ;
        RECT 2891.190 19.920 2891.470 20.200 ;
      LAYER met3 ;
        RECT 2881.000 3009.360 2885.000 3009.960 ;
        RECT 2884.510 3008.810 2884.810 3009.360 ;
        RECT 2891.165 3008.810 2891.495 3008.825 ;
        RECT 2884.510 3008.510 2891.495 3008.810 ;
        RECT 2891.165 3008.495 2891.495 3008.510 ;
        RECT 478.465 20.210 478.795 20.225 ;
        RECT 2891.165 20.210 2891.495 20.225 ;
        RECT 478.465 19.910 2891.495 20.210 ;
        RECT 478.465 19.895 478.795 19.910 ;
        RECT 2891.165 19.895 2891.495 19.910 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.430 15.795 496.710 16.165 ;
        RECT 496.500 2.400 496.640 15.795 ;
        RECT 496.290 -4.800 496.850 2.400 ;
      LAYER via2 ;
        RECT 496.430 15.840 496.710 16.120 ;
      LAYER met3 ;
        RECT 2881.000 3131.080 2885.000 3131.680 ;
        RECT 2884.510 3128.490 2884.810 3131.080 ;
        RECT 2892.750 3128.490 2893.130 3128.500 ;
        RECT 2884.510 3128.190 2893.130 3128.490 ;
        RECT 2892.750 3128.180 2893.130 3128.190 ;
        RECT 496.405 16.130 496.735 16.145 ;
        RECT 2892.750 16.130 2893.130 16.140 ;
        RECT 496.405 15.830 2893.130 16.130 ;
        RECT 496.405 15.815 496.735 15.830 ;
        RECT 2892.750 15.820 2893.130 15.830 ;
      LAYER via3 ;
        RECT 2892.780 3128.180 2893.100 3128.500 ;
        RECT 2892.780 15.820 2893.100 16.140 ;
      LAYER met4 ;
        RECT 2892.775 3128.175 2893.105 3128.505 ;
        RECT 2892.790 16.145 2893.090 3128.175 ;
        RECT 2892.775 15.815 2893.105 16.145 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 513.890 18.600 514.210 18.660 ;
        RECT 2757.770 18.600 2758.090 18.660 ;
        RECT 513.890 18.460 2758.090 18.600 ;
        RECT 513.890 18.400 514.210 18.460 ;
        RECT 2757.770 18.400 2758.090 18.460 ;
      LAYER via ;
        RECT 513.920 18.400 514.180 18.660 ;
        RECT 2757.800 18.400 2758.060 18.660 ;
      LAYER met2 ;
        RECT 2757.830 35.000 2758.110 39.000 ;
        RECT 2757.860 18.690 2758.000 35.000 ;
        RECT 513.920 18.370 514.180 18.690 ;
        RECT 2757.800 18.370 2758.060 18.690 ;
        RECT 513.980 2.400 514.120 18.370 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2620.710 3443.675 2620.990 3444.045 ;
        RECT 2620.780 3435.000 2620.920 3443.675 ;
        RECT 2620.750 3431.000 2621.030 3435.000 ;
        RECT 531.850 37.555 532.130 37.925 ;
        RECT 531.920 2.400 532.060 37.555 ;
        RECT 531.710 -4.800 532.270 2.400 ;
      LAYER via2 ;
        RECT 2620.710 3443.720 2620.990 3444.000 ;
        RECT 531.850 37.600 532.130 37.880 ;
      LAYER met3 ;
        RECT 2620.685 3444.010 2621.015 3444.025 ;
        RECT 2850.430 3444.010 2850.810 3444.020 ;
        RECT 2620.685 3443.710 2850.810 3444.010 ;
        RECT 2620.685 3443.695 2621.015 3443.710 ;
        RECT 2850.430 3443.700 2850.810 3443.710 ;
        RECT 531.825 37.890 532.155 37.905 ;
        RECT 2850.430 37.890 2850.810 37.900 ;
        RECT 531.825 37.590 2850.810 37.890 ;
        RECT 531.825 37.575 532.155 37.590 ;
        RECT 2850.430 37.580 2850.810 37.590 ;
      LAYER via3 ;
        RECT 2850.460 3443.700 2850.780 3444.020 ;
        RECT 2850.460 37.580 2850.780 37.900 ;
      LAYER met4 ;
        RECT 2850.455 3443.695 2850.785 3444.025 ;
        RECT 2850.470 37.905 2850.770 3443.695 ;
        RECT 2850.455 37.575 2850.785 37.905 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2726.510 3444.355 2726.790 3444.725 ;
        RECT 2726.580 3435.000 2726.720 3444.355 ;
        RECT 2726.550 3431.000 2726.830 3435.000 ;
        RECT 549.790 38.235 550.070 38.605 ;
        RECT 549.860 2.400 550.000 38.235 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 2726.510 3444.400 2726.790 3444.680 ;
        RECT 549.790 38.280 550.070 38.560 ;
      LAYER met3 ;
        RECT 2726.485 3444.690 2726.815 3444.705 ;
        RECT 2851.350 3444.690 2851.730 3444.700 ;
        RECT 2726.485 3444.390 2851.730 3444.690 ;
        RECT 2726.485 3444.375 2726.815 3444.390 ;
        RECT 2851.350 3444.380 2851.730 3444.390 ;
        RECT 549.765 38.570 550.095 38.585 ;
        RECT 2851.350 38.570 2851.730 38.580 ;
        RECT 549.765 38.270 2851.730 38.570 ;
        RECT 549.765 38.255 550.095 38.270 ;
        RECT 2851.350 38.260 2851.730 38.270 ;
      LAYER via3 ;
        RECT 2851.380 3444.380 2851.700 3444.700 ;
        RECT 2851.380 38.260 2851.700 38.580 ;
      LAYER met4 ;
        RECT 2851.375 3444.375 2851.705 3444.705 ;
        RECT 2851.390 38.585 2851.690 3444.375 ;
        RECT 2851.375 38.255 2851.705 38.585 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 567.710 19.280 568.030 19.340 ;
        RECT 572.770 19.280 573.090 19.340 ;
        RECT 567.710 19.140 573.090 19.280 ;
        RECT 567.710 19.080 568.030 19.140 ;
        RECT 572.770 19.080 573.090 19.140 ;
      LAYER via ;
        RECT 567.740 19.080 568.000 19.340 ;
        RECT 572.800 19.080 573.060 19.340 ;
      LAYER met2 ;
        RECT 2808.430 35.000 2808.710 39.000 ;
        RECT 2808.460 26.365 2808.600 35.000 ;
        RECT 572.790 25.995 573.070 26.365 ;
        RECT 2808.390 25.995 2808.670 26.365 ;
        RECT 572.860 19.370 573.000 25.995 ;
        RECT 567.740 19.050 568.000 19.370 ;
        RECT 572.800 19.050 573.060 19.370 ;
        RECT 567.800 2.400 567.940 19.050 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 572.790 26.040 573.070 26.320 ;
        RECT 2808.390 26.040 2808.670 26.320 ;
      LAYER met3 ;
        RECT 572.765 26.330 573.095 26.345 ;
        RECT 2808.365 26.330 2808.695 26.345 ;
        RECT 572.765 26.030 2808.695 26.330 ;
        RECT 572.765 26.015 573.095 26.030 ;
        RECT 2808.365 26.015 2808.695 26.030 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 25.830 28.800 26.150 28.860 ;
        RECT 585.650 28.800 585.970 28.860 ;
        RECT 25.830 28.660 585.970 28.800 ;
        RECT 25.830 28.600 26.150 28.660 ;
        RECT 585.650 28.600 585.970 28.660 ;
      LAYER via ;
        RECT 25.860 28.600 26.120 28.860 ;
        RECT 585.680 28.600 585.940 28.860 ;
      LAYER met2 ;
        RECT 25.850 2967.675 26.130 2968.045 ;
        RECT 25.920 28.890 26.060 2967.675 ;
        RECT 25.860 28.570 26.120 28.890 ;
        RECT 585.680 28.570 585.940 28.890 ;
        RECT 585.740 2.400 585.880 28.570 ;
        RECT 585.530 -4.800 586.090 2.400 ;
      LAYER via2 ;
        RECT 25.850 2967.720 26.130 2968.000 ;
      LAYER met3 ;
        RECT 35.000 2970.600 39.000 2971.200 ;
        RECT 25.825 2968.010 26.155 2968.025 ;
        RECT 35.270 2968.010 35.570 2970.600 ;
        RECT 25.825 2967.710 35.570 2968.010 ;
        RECT 25.825 2967.695 26.155 2967.710 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.690 3444.780 45.010 3444.840 ;
        RECT 1987.270 3444.780 1987.590 3444.840 ;
        RECT 44.690 3444.640 1987.590 3444.780 ;
        RECT 44.690 3444.580 45.010 3444.640 ;
        RECT 1987.270 3444.580 1987.590 3444.640 ;
      LAYER via ;
        RECT 44.720 3444.580 44.980 3444.840 ;
        RECT 1987.300 3444.580 1987.560 3444.840 ;
      LAYER met2 ;
        RECT 44.720 3444.550 44.980 3444.870 ;
        RECT 1987.300 3444.550 1987.560 3444.870 ;
        RECT 44.780 17.525 44.920 3444.550 ;
        RECT 1987.360 3435.000 1987.500 3444.550 ;
        RECT 1987.330 3431.000 1987.610 3435.000 ;
        RECT 44.710 17.155 44.990 17.525 ;
        RECT 91.630 17.155 91.910 17.525 ;
        RECT 91.700 2.400 91.840 17.155 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 44.710 17.200 44.990 17.480 ;
        RECT 91.630 17.200 91.910 17.480 ;
      LAYER met3 ;
        RECT 44.685 17.490 45.015 17.505 ;
        RECT 91.605 17.490 91.935 17.505 ;
        RECT 44.685 17.190 91.935 17.490 ;
        RECT 44.685 17.175 45.015 17.190 ;
        RECT 91.605 17.175 91.935 17.190 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.290 18.940 26.610 19.000 ;
        RECT 603.130 18.940 603.450 19.000 ;
        RECT 26.290 18.800 603.450 18.940 ;
        RECT 26.290 18.740 26.610 18.800 ;
        RECT 603.130 18.740 603.450 18.800 ;
      LAYER via ;
        RECT 26.320 18.740 26.580 19.000 ;
        RECT 603.160 18.740 603.420 19.000 ;
      LAYER met2 ;
        RECT 26.310 3070.355 26.590 3070.725 ;
        RECT 26.380 19.030 26.520 3070.355 ;
        RECT 26.320 18.710 26.580 19.030 ;
        RECT 603.160 18.710 603.420 19.030 ;
        RECT 603.220 2.400 603.360 18.710 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 26.310 3070.400 26.590 3070.680 ;
      LAYER met3 ;
        RECT 35.000 3073.280 39.000 3073.880 ;
        RECT 26.285 3070.690 26.615 3070.705 ;
        RECT 35.270 3070.690 35.570 3073.280 ;
        RECT 26.285 3070.390 35.570 3070.690 ;
        RECT 26.285 3070.375 26.615 3070.390 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 621.090 15.115 621.370 15.485 ;
        RECT 621.160 2.400 621.300 15.115 ;
        RECT 620.950 -4.800 621.510 2.400 ;
      LAYER via2 ;
        RECT 621.090 15.160 621.370 15.440 ;
      LAYER met3 ;
        RECT 35.000 3176.640 39.000 3177.240 ;
        RECT 26.950 3174.730 27.330 3174.740 ;
        RECT 35.270 3174.730 35.570 3176.640 ;
        RECT 26.950 3174.430 35.570 3174.730 ;
        RECT 26.950 3174.420 27.330 3174.430 ;
        RECT 26.950 15.450 27.330 15.460 ;
        RECT 621.065 15.450 621.395 15.465 ;
        RECT 26.950 15.150 621.395 15.450 ;
        RECT 26.950 15.140 27.330 15.150 ;
        RECT 621.065 15.135 621.395 15.150 ;
      LAYER via3 ;
        RECT 26.980 3174.420 27.300 3174.740 ;
        RECT 26.980 15.140 27.300 15.460 ;
      LAYER met4 ;
        RECT 26.975 3174.415 27.305 3174.745 ;
        RECT 26.990 15.465 27.290 3174.415 ;
        RECT 26.975 15.135 27.305 15.465 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 46.530 3444.440 46.850 3444.500 ;
        RECT 2093.070 3444.440 2093.390 3444.500 ;
        RECT 46.530 3444.300 2093.390 3444.440 ;
        RECT 46.530 3444.240 46.850 3444.300 ;
        RECT 2093.070 3444.240 2093.390 3444.300 ;
      LAYER via ;
        RECT 46.560 3444.240 46.820 3444.500 ;
        RECT 2093.100 3444.240 2093.360 3444.500 ;
      LAYER met2 ;
        RECT 46.560 3444.210 46.820 3444.530 ;
        RECT 2093.100 3444.210 2093.360 3444.530 ;
        RECT 46.620 18.205 46.760 3444.210 ;
        RECT 2093.160 3435.000 2093.300 3444.210 ;
        RECT 2093.130 3431.000 2093.410 3435.000 ;
        RECT 46.550 17.835 46.830 18.205 ;
        RECT 115.550 17.835 115.830 18.205 ;
        RECT 115.620 2.400 115.760 17.835 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 46.550 17.880 46.830 18.160 ;
        RECT 115.550 17.880 115.830 18.160 ;
      LAYER met3 ;
        RECT 46.525 18.170 46.855 18.185 ;
        RECT 115.525 18.170 115.855 18.185 ;
        RECT 46.525 17.870 115.855 18.170 ;
        RECT 46.525 17.855 46.855 17.870 ;
        RECT 115.525 17.855 115.855 17.870 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 139.450 17.240 139.770 17.300 ;
        RECT 2894.850 17.240 2895.170 17.300 ;
        RECT 139.450 17.100 2895.170 17.240 ;
        RECT 139.450 17.040 139.770 17.100 ;
        RECT 2894.850 17.040 2895.170 17.100 ;
      LAYER via ;
        RECT 139.480 17.040 139.740 17.300 ;
        RECT 2894.880 17.040 2895.140 17.300 ;
      LAYER met2 ;
        RECT 2894.870 2035.395 2895.150 2035.765 ;
        RECT 2894.940 17.330 2895.080 2035.395 ;
        RECT 139.480 17.010 139.740 17.330 ;
        RECT 2894.880 17.010 2895.140 17.330 ;
        RECT 139.540 2.400 139.680 17.010 ;
        RECT 139.330 -4.800 139.890 2.400 ;
      LAYER via2 ;
        RECT 2894.870 2035.440 2895.150 2035.720 ;
      LAYER met3 ;
        RECT 2881.000 2038.320 2885.000 2038.920 ;
        RECT 2884.510 2035.730 2884.810 2038.320 ;
        RECT 2894.845 2035.730 2895.175 2035.745 ;
        RECT 2884.510 2035.430 2895.175 2035.730 ;
        RECT 2894.845 2035.415 2895.175 2035.430 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 157.390 17.580 157.710 17.640 ;
        RECT 2894.390 17.580 2894.710 17.640 ;
        RECT 157.390 17.440 2894.710 17.580 ;
        RECT 157.390 17.380 157.710 17.440 ;
        RECT 2894.390 17.380 2894.710 17.440 ;
      LAYER via ;
        RECT 157.420 17.380 157.680 17.640 ;
        RECT 2894.420 17.380 2894.680 17.640 ;
      LAYER met2 ;
        RECT 2894.410 2156.435 2894.690 2156.805 ;
        RECT 2894.480 17.670 2894.620 2156.435 ;
        RECT 157.420 17.350 157.680 17.670 ;
        RECT 2894.420 17.350 2894.680 17.670 ;
        RECT 157.480 2.400 157.620 17.350 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 2894.410 2156.480 2894.690 2156.760 ;
      LAYER met3 ;
        RECT 2881.000 2159.360 2885.000 2159.960 ;
        RECT 2884.510 2156.770 2884.810 2159.360 ;
        RECT 2894.385 2156.770 2894.715 2156.785 ;
        RECT 2884.510 2156.470 2894.715 2156.770 ;
        RECT 2894.385 2156.455 2894.715 2156.470 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2605.110 35.000 2605.390 39.000 ;
        RECT 2605.140 25.685 2605.280 35.000 ;
        RECT 174.890 25.315 175.170 25.685 ;
        RECT 2605.070 25.315 2605.350 25.685 ;
        RECT 174.960 2.400 175.100 25.315 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 174.890 25.360 175.170 25.640 ;
        RECT 2605.070 25.360 2605.350 25.640 ;
      LAYER met3 ;
        RECT 174.865 25.650 175.195 25.665 ;
        RECT 2605.045 25.650 2605.375 25.665 ;
        RECT 174.865 25.350 2605.375 25.650 ;
        RECT 174.865 25.335 175.195 25.350 ;
        RECT 2605.045 25.335 2605.375 25.350 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2655.710 35.000 2655.990 39.000 ;
        RECT 2655.740 25.005 2655.880 35.000 ;
        RECT 192.830 24.635 193.110 25.005 ;
        RECT 2655.670 24.635 2655.950 25.005 ;
        RECT 192.900 2.400 193.040 24.635 ;
        RECT 192.690 -4.800 193.250 2.400 ;
      LAYER via2 ;
        RECT 192.830 24.680 193.110 24.960 ;
        RECT 2655.670 24.680 2655.950 24.960 ;
      LAYER met3 ;
        RECT 192.805 24.970 193.135 24.985 ;
        RECT 2655.645 24.970 2655.975 24.985 ;
        RECT 192.805 24.670 2655.975 24.970 ;
        RECT 192.805 24.655 193.135 24.670 ;
        RECT 2655.645 24.655 2655.975 24.670 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2893.950 2278.155 2894.230 2278.525 ;
        RECT 2894.020 18.885 2894.160 2278.155 ;
        RECT 210.770 18.515 211.050 18.885 ;
        RECT 2893.950 18.515 2894.230 18.885 ;
        RECT 210.840 2.400 210.980 18.515 ;
        RECT 210.630 -4.800 211.190 2.400 ;
      LAYER via2 ;
        RECT 2893.950 2278.200 2894.230 2278.480 ;
        RECT 210.770 18.560 211.050 18.840 ;
        RECT 2893.950 18.560 2894.230 18.840 ;
      LAYER met3 ;
        RECT 2881.000 2281.080 2885.000 2281.680 ;
        RECT 2884.510 2278.490 2884.810 2281.080 ;
        RECT 2893.925 2278.490 2894.255 2278.505 ;
        RECT 2884.510 2278.190 2894.255 2278.490 ;
        RECT 2893.925 2278.175 2894.255 2278.190 ;
        RECT 210.745 18.850 211.075 18.865 ;
        RECT 2893.925 18.850 2894.255 18.865 ;
        RECT 210.745 18.550 2894.255 18.850 ;
        RECT 210.745 18.535 211.075 18.550 ;
        RECT 2893.925 18.535 2894.255 18.550 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 25.370 15.880 25.690 15.940 ;
        RECT 228.690 15.880 229.010 15.940 ;
        RECT 25.370 15.740 229.010 15.880 ;
        RECT 25.370 15.680 25.690 15.740 ;
        RECT 228.690 15.680 229.010 15.740 ;
      LAYER via ;
        RECT 25.400 15.680 25.660 15.940 ;
        RECT 228.720 15.680 228.980 15.940 ;
      LAYER met2 ;
        RECT 25.390 2555.595 25.670 2555.965 ;
        RECT 25.460 15.970 25.600 2555.595 ;
        RECT 25.400 15.650 25.660 15.970 ;
        RECT 228.720 15.650 228.980 15.970 ;
        RECT 228.780 2.400 228.920 15.650 ;
        RECT 228.570 -4.800 229.130 2.400 ;
      LAYER via2 ;
        RECT 25.390 2555.640 25.670 2555.920 ;
      LAYER met3 ;
        RECT 35.000 2558.520 39.000 2559.120 ;
        RECT 25.365 2555.930 25.695 2555.945 ;
        RECT 35.270 2555.930 35.570 2558.520 ;
        RECT 25.365 2555.630 35.570 2555.930 ;
        RECT 25.365 2555.615 25.695 2555.630 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 50.210 18.600 50.530 18.660 ;
        RECT 465.590 18.600 465.910 18.660 ;
        RECT 50.210 18.460 465.910 18.600 ;
        RECT 50.210 18.400 50.530 18.460 ;
        RECT 465.590 18.400 465.910 18.460 ;
      LAYER via ;
        RECT 50.240 18.400 50.500 18.660 ;
        RECT 465.620 18.400 465.880 18.660 ;
      LAYER met2 ;
        RECT 467.490 35.770 467.770 39.000 ;
        RECT 465.680 35.630 467.770 35.770 ;
        RECT 465.680 18.690 465.820 35.630 ;
        RECT 467.490 35.000 467.770 35.630 ;
        RECT 50.240 18.370 50.500 18.690 ;
        RECT 465.620 18.370 465.880 18.690 ;
        RECT 50.300 2.400 50.440 18.370 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 252.610 14.860 252.930 14.920 ;
        RECT 976.190 14.860 976.510 14.920 ;
        RECT 252.610 14.720 976.510 14.860 ;
        RECT 252.610 14.660 252.930 14.720 ;
        RECT 976.190 14.660 976.510 14.720 ;
      LAYER via ;
        RECT 252.640 14.660 252.900 14.920 ;
        RECT 976.220 14.660 976.480 14.920 ;
      LAYER met2 ;
        RECT 976.250 35.000 976.530 39.000 ;
        RECT 976.280 14.950 976.420 35.000 ;
        RECT 252.640 14.630 252.900 14.950 ;
        RECT 976.220 14.630 976.480 14.950 ;
        RECT 252.700 2.400 252.840 14.630 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 513.045 16.745 513.215 19.635 ;
      LAYER mcon ;
        RECT 513.045 19.465 513.215 19.635 ;
      LAYER met1 ;
        RECT 552.070 20.980 552.390 21.040 ;
        RECT 1027.250 20.980 1027.570 21.040 ;
        RECT 552.070 20.840 1027.570 20.980 ;
        RECT 552.070 20.780 552.390 20.840 ;
        RECT 1027.250 20.780 1027.570 20.840 ;
        RECT 512.985 19.620 513.275 19.665 ;
        RECT 552.070 19.620 552.390 19.680 ;
        RECT 512.985 19.480 552.390 19.620 ;
        RECT 512.985 19.435 513.275 19.480 ;
        RECT 552.070 19.420 552.390 19.480 ;
        RECT 270.090 16.900 270.410 16.960 ;
        RECT 512.985 16.900 513.275 16.945 ;
        RECT 270.090 16.760 513.275 16.900 ;
        RECT 270.090 16.700 270.410 16.760 ;
        RECT 512.985 16.715 513.275 16.760 ;
      LAYER via ;
        RECT 552.100 20.780 552.360 21.040 ;
        RECT 1027.280 20.780 1027.540 21.040 ;
        RECT 552.100 19.420 552.360 19.680 ;
        RECT 270.120 16.700 270.380 16.960 ;
      LAYER met2 ;
        RECT 1027.310 35.000 1027.590 39.000 ;
        RECT 1027.340 21.070 1027.480 35.000 ;
        RECT 552.100 20.750 552.360 21.070 ;
        RECT 1027.280 20.750 1027.540 21.070 ;
        RECT 552.160 19.710 552.300 20.750 ;
        RECT 552.100 19.390 552.360 19.710 ;
        RECT 270.120 16.670 270.380 16.990 ;
        RECT 270.180 2.400 270.320 16.670 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.030 15.200 288.350 15.260 ;
        RECT 1077.850 15.200 1078.170 15.260 ;
        RECT 288.030 15.060 1078.170 15.200 ;
        RECT 288.030 15.000 288.350 15.060 ;
        RECT 1077.850 15.000 1078.170 15.060 ;
      LAYER via ;
        RECT 288.060 15.000 288.320 15.260 ;
        RECT 1077.880 15.000 1078.140 15.260 ;
      LAYER met2 ;
        RECT 1077.910 35.000 1078.190 39.000 ;
        RECT 1077.940 15.290 1078.080 35.000 ;
        RECT 288.060 14.970 288.320 15.290 ;
        RECT 1077.880 14.970 1078.140 15.290 ;
        RECT 288.120 2.400 288.260 14.970 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 348.825 16.065 348.995 20.315 ;
      LAYER mcon ;
        RECT 348.825 20.145 348.995 20.315 ;
      LAYER met1 ;
        RECT 569.550 22.000 569.870 22.060 ;
        RECT 1128.910 22.000 1129.230 22.060 ;
        RECT 569.550 21.860 1129.230 22.000 ;
        RECT 569.550 21.800 569.870 21.860 ;
        RECT 1128.910 21.800 1129.230 21.860 ;
        RECT 348.765 20.300 349.055 20.345 ;
        RECT 569.550 20.300 569.870 20.360 ;
        RECT 348.765 20.160 569.870 20.300 ;
        RECT 348.765 20.115 349.055 20.160 ;
        RECT 569.550 20.100 569.870 20.160 ;
        RECT 305.970 16.560 306.290 16.620 ;
        RECT 305.970 16.420 348.060 16.560 ;
        RECT 305.970 16.360 306.290 16.420 ;
        RECT 347.920 16.220 348.060 16.420 ;
        RECT 348.765 16.220 349.055 16.265 ;
        RECT 347.920 16.080 349.055 16.220 ;
        RECT 348.765 16.035 349.055 16.080 ;
      LAYER via ;
        RECT 569.580 21.800 569.840 22.060 ;
        RECT 1128.940 21.800 1129.200 22.060 ;
        RECT 569.580 20.100 569.840 20.360 ;
        RECT 306.000 16.360 306.260 16.620 ;
      LAYER met2 ;
        RECT 1128.970 35.000 1129.250 39.000 ;
        RECT 1129.000 22.090 1129.140 35.000 ;
        RECT 569.580 21.770 569.840 22.090 ;
        RECT 1128.940 21.770 1129.200 22.090 ;
        RECT 569.640 20.390 569.780 21.770 ;
        RECT 569.580 20.070 569.840 20.390 ;
        RECT 306.000 16.330 306.260 16.650 ;
        RECT 306.060 2.400 306.200 16.330 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 15.540 324.230 15.600 ;
        RECT 1179.970 15.540 1180.290 15.600 ;
        RECT 323.910 15.400 1180.290 15.540 ;
        RECT 323.910 15.340 324.230 15.400 ;
        RECT 1179.970 15.340 1180.290 15.400 ;
      LAYER via ;
        RECT 323.940 15.340 324.200 15.600 ;
        RECT 1180.000 15.340 1180.260 15.600 ;
      LAYER met2 ;
        RECT 1180.030 35.000 1180.310 39.000 ;
        RECT 1180.060 15.630 1180.200 35.000 ;
        RECT 323.940 15.310 324.200 15.630 ;
        RECT 1180.000 15.310 1180.260 15.630 ;
        RECT 324.000 2.400 324.140 15.310 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 23.020 341.710 23.080 ;
        RECT 1230.570 23.020 1230.890 23.080 ;
        RECT 341.390 22.880 1230.890 23.020 ;
        RECT 341.390 22.820 341.710 22.880 ;
        RECT 1230.570 22.820 1230.890 22.880 ;
      LAYER via ;
        RECT 341.420 22.820 341.680 23.080 ;
        RECT 1230.600 22.820 1230.860 23.080 ;
      LAYER met2 ;
        RECT 1230.630 35.000 1230.910 39.000 ;
        RECT 1230.660 23.110 1230.800 35.000 ;
        RECT 341.420 22.790 341.680 23.110 ;
        RECT 1230.600 22.790 1230.860 23.110 ;
        RECT 341.480 2.400 341.620 22.790 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 359.330 15.880 359.650 15.940 ;
        RECT 1281.630 15.880 1281.950 15.940 ;
        RECT 359.330 15.740 1281.950 15.880 ;
        RECT 359.330 15.680 359.650 15.740 ;
        RECT 1281.630 15.680 1281.950 15.740 ;
      LAYER via ;
        RECT 359.360 15.680 359.620 15.940 ;
        RECT 1281.660 15.680 1281.920 15.940 ;
      LAYER met2 ;
        RECT 1281.690 35.000 1281.970 39.000 ;
        RECT 1281.720 15.970 1281.860 35.000 ;
        RECT 359.360 15.650 359.620 15.970 ;
        RECT 1281.660 15.650 1281.920 15.970 ;
        RECT 359.420 2.400 359.560 15.650 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 377.270 23.360 377.590 23.420 ;
        RECT 1332.690 23.360 1333.010 23.420 ;
        RECT 377.270 23.220 1333.010 23.360 ;
        RECT 377.270 23.160 377.590 23.220 ;
        RECT 1332.690 23.160 1333.010 23.220 ;
      LAYER via ;
        RECT 377.300 23.160 377.560 23.420 ;
        RECT 1332.720 23.160 1332.980 23.420 ;
      LAYER met2 ;
        RECT 1332.750 35.000 1333.030 39.000 ;
        RECT 1332.780 23.450 1332.920 35.000 ;
        RECT 377.300 23.130 377.560 23.450 ;
        RECT 1332.720 23.130 1332.980 23.450 ;
        RECT 377.360 2.400 377.500 23.130 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 395.210 16.220 395.530 16.280 ;
        RECT 1383.290 16.220 1383.610 16.280 ;
        RECT 395.210 16.080 1383.610 16.220 ;
        RECT 395.210 16.020 395.530 16.080 ;
        RECT 1383.290 16.020 1383.610 16.080 ;
      LAYER via ;
        RECT 395.240 16.020 395.500 16.280 ;
        RECT 1383.320 16.020 1383.580 16.280 ;
      LAYER met2 ;
        RECT 1383.350 35.000 1383.630 39.000 ;
        RECT 1383.380 16.310 1383.520 35.000 ;
        RECT 395.240 15.990 395.500 16.310 ;
        RECT 1383.320 15.990 1383.580 16.310 ;
        RECT 395.300 2.400 395.440 15.990 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 413.150 23.700 413.470 23.760 ;
        RECT 1434.350 23.700 1434.670 23.760 ;
        RECT 413.150 23.560 1434.670 23.700 ;
        RECT 413.150 23.500 413.470 23.560 ;
        RECT 1434.350 23.500 1434.670 23.560 ;
      LAYER via ;
        RECT 413.180 23.500 413.440 23.760 ;
        RECT 1434.380 23.500 1434.640 23.760 ;
      LAYER met2 ;
        RECT 1434.410 35.000 1434.690 39.000 ;
        RECT 1434.440 23.790 1434.580 35.000 ;
        RECT 413.180 23.470 413.440 23.790 ;
        RECT 1434.380 23.470 1434.640 23.790 ;
        RECT 413.240 2.400 413.380 23.470 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 82.945 17.425 83.115 19.295 ;
        RECT 130.785 17.425 130.955 19.295 ;
        RECT 179.545 14.365 179.715 19.295 ;
        RECT 227.385 14.705 227.555 19.295 ;
        RECT 276.145 15.725 276.315 19.295 ;
        RECT 323.985 16.065 324.155 19.295 ;
        RECT 372.745 19.125 372.915 20.655 ;
        RECT 420.585 19.125 420.755 20.655 ;
        RECT 512.585 19.465 512.755 20.995 ;
      LAYER mcon ;
        RECT 512.585 20.825 512.755 20.995 ;
        RECT 372.745 20.485 372.915 20.655 ;
        RECT 82.945 19.125 83.115 19.295 ;
        RECT 130.785 19.125 130.955 19.295 ;
        RECT 179.545 19.125 179.715 19.295 ;
        RECT 227.385 19.125 227.555 19.295 ;
        RECT 276.145 19.125 276.315 19.295 ;
        RECT 323.985 19.125 324.155 19.295 ;
        RECT 420.585 20.485 420.755 20.655 ;
      LAYER met1 ;
        RECT 512.525 20.980 512.815 21.025 ;
        RECT 518.030 20.980 518.350 21.040 ;
        RECT 512.525 20.840 518.350 20.980 ;
        RECT 512.525 20.795 512.815 20.840 ;
        RECT 518.030 20.780 518.350 20.840 ;
        RECT 372.685 20.640 372.975 20.685 ;
        RECT 420.525 20.640 420.815 20.685 ;
        RECT 372.685 20.500 420.815 20.640 ;
        RECT 372.685 20.455 372.975 20.500 ;
        RECT 420.525 20.455 420.815 20.500 ;
        RECT 512.525 19.620 512.815 19.665 ;
        RECT 493.280 19.480 512.815 19.620 ;
        RECT 74.130 19.280 74.450 19.340 ;
        RECT 82.885 19.280 83.175 19.325 ;
        RECT 74.130 19.140 83.175 19.280 ;
        RECT 74.130 19.080 74.450 19.140 ;
        RECT 82.885 19.095 83.175 19.140 ;
        RECT 130.725 19.280 131.015 19.325 ;
        RECT 179.485 19.280 179.775 19.325 ;
        RECT 130.725 19.140 179.775 19.280 ;
        RECT 130.725 19.095 131.015 19.140 ;
        RECT 179.485 19.095 179.775 19.140 ;
        RECT 227.325 19.280 227.615 19.325 ;
        RECT 276.085 19.280 276.375 19.325 ;
        RECT 227.325 19.140 276.375 19.280 ;
        RECT 227.325 19.095 227.615 19.140 ;
        RECT 276.085 19.095 276.375 19.140 ;
        RECT 323.925 19.280 324.215 19.325 ;
        RECT 372.685 19.280 372.975 19.325 ;
        RECT 323.925 19.140 372.975 19.280 ;
        RECT 323.925 19.095 324.215 19.140 ;
        RECT 372.685 19.095 372.975 19.140 ;
        RECT 420.525 19.280 420.815 19.325 ;
        RECT 493.280 19.280 493.420 19.480 ;
        RECT 512.525 19.435 512.815 19.480 ;
        RECT 420.525 19.140 493.420 19.280 ;
        RECT 420.525 19.095 420.815 19.140 ;
        RECT 82.885 17.580 83.175 17.625 ;
        RECT 130.725 17.580 131.015 17.625 ;
        RECT 82.885 17.440 131.015 17.580 ;
        RECT 82.885 17.395 83.175 17.440 ;
        RECT 130.725 17.395 131.015 17.440 ;
        RECT 323.925 16.035 324.215 16.265 ;
        RECT 276.085 15.880 276.375 15.925 ;
        RECT 324.000 15.880 324.140 16.035 ;
        RECT 276.085 15.740 324.140 15.880 ;
        RECT 276.085 15.695 276.375 15.740 ;
        RECT 227.325 14.860 227.615 14.905 ;
        RECT 187.380 14.720 227.615 14.860 ;
        RECT 179.485 14.520 179.775 14.565 ;
        RECT 187.380 14.520 187.520 14.720 ;
        RECT 227.325 14.675 227.615 14.720 ;
        RECT 179.485 14.380 187.520 14.520 ;
        RECT 179.485 14.335 179.775 14.380 ;
      LAYER via ;
        RECT 518.060 20.780 518.320 21.040 ;
        RECT 74.160 19.080 74.420 19.340 ;
      LAYER met2 ;
        RECT 518.090 35.000 518.370 39.000 ;
        RECT 518.120 21.070 518.260 35.000 ;
        RECT 518.060 20.750 518.320 21.070 ;
        RECT 74.160 19.050 74.420 19.370 ;
        RECT 74.220 2.400 74.360 19.050 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 430.630 16.560 430.950 16.620 ;
        RECT 1485.410 16.560 1485.730 16.620 ;
        RECT 430.630 16.420 1485.730 16.560 ;
        RECT 430.630 16.360 430.950 16.420 ;
        RECT 1485.410 16.360 1485.730 16.420 ;
      LAYER via ;
        RECT 430.660 16.360 430.920 16.620 ;
        RECT 1485.440 16.360 1485.700 16.620 ;
      LAYER met2 ;
        RECT 1485.470 35.000 1485.750 39.000 ;
        RECT 1485.500 16.650 1485.640 35.000 ;
        RECT 430.660 16.330 430.920 16.650 ;
        RECT 1485.440 16.330 1485.700 16.650 ;
        RECT 430.720 2.400 430.860 16.330 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.570 27.440 448.890 27.500 ;
        RECT 1536.010 27.440 1536.330 27.500 ;
        RECT 448.570 27.300 1536.330 27.440 ;
        RECT 448.570 27.240 448.890 27.300 ;
        RECT 1536.010 27.240 1536.330 27.300 ;
      LAYER via ;
        RECT 448.600 27.240 448.860 27.500 ;
        RECT 1536.040 27.240 1536.300 27.500 ;
      LAYER met2 ;
        RECT 1536.070 35.000 1536.350 39.000 ;
        RECT 1536.100 27.530 1536.240 35.000 ;
        RECT 448.600 27.210 448.860 27.530 ;
        RECT 1536.040 27.210 1536.300 27.530 ;
        RECT 448.660 2.400 448.800 27.210 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 513.505 16.745 513.675 18.615 ;
      LAYER mcon ;
        RECT 513.505 18.445 513.675 18.615 ;
      LAYER met1 ;
        RECT 466.510 18.600 466.830 18.660 ;
        RECT 513.445 18.600 513.735 18.645 ;
        RECT 466.510 18.460 513.735 18.600 ;
        RECT 466.510 18.400 466.830 18.460 ;
        RECT 513.445 18.415 513.735 18.460 ;
        RECT 513.445 16.900 513.735 16.945 ;
        RECT 1587.070 16.900 1587.390 16.960 ;
        RECT 513.445 16.760 1587.390 16.900 ;
        RECT 513.445 16.715 513.735 16.760 ;
        RECT 1587.070 16.700 1587.390 16.760 ;
      LAYER via ;
        RECT 466.540 18.400 466.800 18.660 ;
        RECT 1587.100 16.700 1587.360 16.960 ;
      LAYER met2 ;
        RECT 1587.130 35.000 1587.410 39.000 ;
        RECT 466.540 18.370 466.800 18.690 ;
        RECT 466.600 2.400 466.740 18.370 ;
        RECT 1587.160 16.990 1587.300 35.000 ;
        RECT 1587.100 16.670 1587.360 16.990 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 484.450 27.100 484.770 27.160 ;
        RECT 1637.670 27.100 1637.990 27.160 ;
        RECT 484.450 26.960 1637.990 27.100 ;
        RECT 484.450 26.900 484.770 26.960 ;
        RECT 1637.670 26.900 1637.990 26.960 ;
      LAYER via ;
        RECT 484.480 26.900 484.740 27.160 ;
        RECT 1637.700 26.900 1637.960 27.160 ;
      LAYER met2 ;
        RECT 1637.730 35.000 1638.010 39.000 ;
        RECT 1637.760 27.190 1637.900 35.000 ;
        RECT 484.480 26.870 484.740 27.190 ;
        RECT 1637.700 26.870 1637.960 27.190 ;
        RECT 484.540 2.400 484.680 26.870 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 502.390 20.640 502.710 20.700 ;
        RECT 1688.730 20.640 1689.050 20.700 ;
        RECT 502.390 20.500 1689.050 20.640 ;
        RECT 502.390 20.440 502.710 20.500 ;
        RECT 1688.730 20.440 1689.050 20.500 ;
      LAYER via ;
        RECT 502.420 20.440 502.680 20.700 ;
        RECT 1688.760 20.440 1689.020 20.700 ;
      LAYER met2 ;
        RECT 1688.790 35.000 1689.070 39.000 ;
        RECT 1688.820 20.730 1688.960 35.000 ;
        RECT 502.420 20.410 502.680 20.730 ;
        RECT 1688.760 20.410 1689.020 20.730 ;
        RECT 502.480 2.400 502.620 20.410 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 519.870 26.760 520.190 26.820 ;
        RECT 1739.790 26.760 1740.110 26.820 ;
        RECT 519.870 26.620 1740.110 26.760 ;
        RECT 519.870 26.560 520.190 26.620 ;
        RECT 1739.790 26.560 1740.110 26.620 ;
      LAYER via ;
        RECT 519.900 26.560 520.160 26.820 ;
        RECT 1739.820 26.560 1740.080 26.820 ;
      LAYER met2 ;
        RECT 1739.850 35.000 1740.130 39.000 ;
        RECT 1739.880 26.850 1740.020 35.000 ;
        RECT 519.900 26.530 520.160 26.850 ;
        RECT 1739.820 26.530 1740.080 26.850 ;
        RECT 519.960 2.400 520.100 26.530 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1790.390 20.300 1790.710 20.360 ;
        RECT 589.420 20.160 1790.710 20.300 ;
        RECT 537.810 19.960 538.130 20.020 ;
        RECT 589.420 19.960 589.560 20.160 ;
        RECT 1790.390 20.100 1790.710 20.160 ;
        RECT 537.810 19.820 589.560 19.960 ;
        RECT 537.810 19.760 538.130 19.820 ;
      LAYER via ;
        RECT 537.840 19.760 538.100 20.020 ;
        RECT 1790.420 20.100 1790.680 20.360 ;
      LAYER met2 ;
        RECT 1790.450 35.000 1790.730 39.000 ;
        RECT 1790.480 20.390 1790.620 35.000 ;
        RECT 1790.420 20.070 1790.680 20.390 ;
        RECT 537.840 19.730 538.100 20.050 ;
        RECT 537.900 2.400 538.040 19.730 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1841.450 19.960 1841.770 20.020 ;
        RECT 589.880 19.820 1841.770 19.960 ;
        RECT 555.750 19.620 556.070 19.680 ;
        RECT 589.880 19.620 590.020 19.820 ;
        RECT 1841.450 19.760 1841.770 19.820 ;
        RECT 555.750 19.480 590.020 19.620 ;
        RECT 555.750 19.420 556.070 19.480 ;
      LAYER via ;
        RECT 555.780 19.420 556.040 19.680 ;
        RECT 1841.480 19.760 1841.740 20.020 ;
      LAYER met2 ;
        RECT 1841.510 35.000 1841.790 39.000 ;
        RECT 1841.540 20.050 1841.680 35.000 ;
        RECT 1841.480 19.730 1841.740 20.050 ;
        RECT 555.780 19.390 556.040 19.710 ;
        RECT 555.840 2.400 555.980 19.390 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1892.510 19.620 1892.830 19.680 ;
        RECT 590.340 19.480 1892.830 19.620 ;
        RECT 573.690 19.280 574.010 19.340 ;
        RECT 590.340 19.280 590.480 19.480 ;
        RECT 1892.510 19.420 1892.830 19.480 ;
        RECT 573.690 19.140 590.480 19.280 ;
        RECT 573.690 19.080 574.010 19.140 ;
      LAYER via ;
        RECT 573.720 19.080 573.980 19.340 ;
        RECT 1892.540 19.420 1892.800 19.680 ;
      LAYER met2 ;
        RECT 1892.570 35.000 1892.850 39.000 ;
        RECT 1892.600 19.710 1892.740 35.000 ;
        RECT 1892.540 19.390 1892.800 19.710 ;
        RECT 573.720 19.050 573.980 19.370 ;
        RECT 573.780 2.400 573.920 19.050 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 591.170 19.280 591.490 19.340 ;
        RECT 1943.110 19.280 1943.430 19.340 ;
        RECT 591.170 19.140 1943.430 19.280 ;
        RECT 591.170 19.080 591.490 19.140 ;
        RECT 1943.110 19.080 1943.430 19.140 ;
      LAYER via ;
        RECT 591.200 19.080 591.460 19.340 ;
        RECT 1943.140 19.080 1943.400 19.340 ;
      LAYER met2 ;
        RECT 1943.170 35.000 1943.450 39.000 ;
        RECT 1943.200 19.370 1943.340 35.000 ;
        RECT 591.200 19.050 591.460 19.370 ;
        RECT 1943.140 19.050 1943.400 19.370 ;
        RECT 591.260 2.400 591.400 19.050 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 97.590 22.000 97.910 22.060 ;
        RECT 565.410 22.000 565.730 22.060 ;
        RECT 97.590 21.860 565.730 22.000 ;
        RECT 97.590 21.800 97.910 21.860 ;
        RECT 565.410 21.800 565.730 21.860 ;
      LAYER via ;
        RECT 97.620 21.800 97.880 22.060 ;
        RECT 565.440 21.800 565.700 22.060 ;
      LAYER met2 ;
        RECT 569.150 35.770 569.430 39.000 ;
        RECT 565.960 35.630 569.430 35.770 ;
        RECT 565.960 22.850 566.100 35.630 ;
        RECT 569.150 35.000 569.430 35.630 ;
        RECT 565.500 22.710 566.100 22.850 ;
        RECT 565.500 22.090 565.640 22.710 ;
        RECT 97.620 21.770 97.880 22.090 ;
        RECT 565.440 21.770 565.700 22.090 ;
        RECT 97.680 2.400 97.820 21.770 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 620.610 26.420 620.930 26.480 ;
        RECT 1994.170 26.420 1994.490 26.480 ;
        RECT 620.610 26.280 1994.490 26.420 ;
        RECT 620.610 26.220 620.930 26.280 ;
        RECT 1994.170 26.220 1994.490 26.280 ;
        RECT 609.110 18.940 609.430 19.000 ;
        RECT 620.610 18.940 620.930 19.000 ;
        RECT 609.110 18.800 620.930 18.940 ;
        RECT 609.110 18.740 609.430 18.800 ;
        RECT 620.610 18.740 620.930 18.800 ;
      LAYER via ;
        RECT 620.640 26.220 620.900 26.480 ;
        RECT 1994.200 26.220 1994.460 26.480 ;
        RECT 609.140 18.740 609.400 19.000 ;
        RECT 620.640 18.740 620.900 19.000 ;
      LAYER met2 ;
        RECT 1994.230 35.000 1994.510 39.000 ;
        RECT 1994.260 26.510 1994.400 35.000 ;
        RECT 620.640 26.190 620.900 26.510 ;
        RECT 1994.200 26.190 1994.460 26.510 ;
        RECT 620.700 19.030 620.840 26.190 ;
        RECT 609.140 18.710 609.400 19.030 ;
        RECT 620.640 18.710 620.900 19.030 ;
        RECT 609.200 2.400 609.340 18.710 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.050 18.940 627.370 19.000 ;
        RECT 2045.230 18.940 2045.550 19.000 ;
        RECT 627.050 18.800 2045.550 18.940 ;
        RECT 627.050 18.740 627.370 18.800 ;
        RECT 2045.230 18.740 2045.550 18.800 ;
      LAYER via ;
        RECT 627.080 18.740 627.340 19.000 ;
        RECT 2045.260 18.740 2045.520 19.000 ;
      LAYER met2 ;
        RECT 2045.290 35.000 2045.570 39.000 ;
        RECT 2045.320 19.030 2045.460 35.000 ;
        RECT 627.080 18.710 627.340 19.030 ;
        RECT 2045.260 18.710 2045.520 19.030 ;
        RECT 627.140 2.400 627.280 18.710 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 26.420 121.830 26.480 ;
        RECT 620.150 26.420 620.470 26.480 ;
        RECT 121.510 26.280 620.470 26.420 ;
        RECT 121.510 26.220 121.830 26.280 ;
        RECT 620.150 26.220 620.470 26.280 ;
      LAYER via ;
        RECT 121.540 26.220 121.800 26.480 ;
        RECT 620.180 26.220 620.440 26.480 ;
      LAYER met2 ;
        RECT 620.210 35.000 620.490 39.000 ;
        RECT 620.240 26.510 620.380 35.000 ;
        RECT 121.540 26.190 121.800 26.510 ;
        RECT 620.180 26.190 620.440 26.510 ;
        RECT 121.600 2.400 121.740 26.190 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 145.430 21.320 145.750 21.380 ;
        RECT 670.750 21.320 671.070 21.380 ;
        RECT 145.430 21.180 671.070 21.320 ;
        RECT 145.430 21.120 145.750 21.180 ;
        RECT 670.750 21.120 671.070 21.180 ;
      LAYER via ;
        RECT 145.460 21.120 145.720 21.380 ;
        RECT 670.780 21.120 671.040 21.380 ;
      LAYER met2 ;
        RECT 670.810 35.000 671.090 39.000 ;
        RECT 670.840 21.410 670.980 35.000 ;
        RECT 145.460 21.090 145.720 21.410 ;
        RECT 670.780 21.090 671.040 21.410 ;
        RECT 145.520 2.400 145.660 21.090 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 163.370 21.660 163.690 21.720 ;
        RECT 721.810 21.660 722.130 21.720 ;
        RECT 163.370 21.520 722.130 21.660 ;
        RECT 163.370 21.460 163.690 21.520 ;
        RECT 721.810 21.460 722.130 21.520 ;
      LAYER via ;
        RECT 163.400 21.460 163.660 21.720 ;
        RECT 721.840 21.460 722.100 21.720 ;
      LAYER met2 ;
        RECT 721.870 35.000 722.150 39.000 ;
        RECT 721.900 21.750 722.040 35.000 ;
        RECT 163.400 21.430 163.660 21.750 ;
        RECT 721.840 21.430 722.100 21.750 ;
        RECT 163.460 2.400 163.600 21.430 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 180.850 14.180 181.170 14.240 ;
        RECT 772.870 14.180 773.190 14.240 ;
        RECT 180.850 14.040 773.190 14.180 ;
        RECT 180.850 13.980 181.170 14.040 ;
        RECT 772.870 13.980 773.190 14.040 ;
      LAYER via ;
        RECT 180.880 13.980 181.140 14.240 ;
        RECT 772.900 13.980 773.160 14.240 ;
      LAYER met2 ;
        RECT 772.930 35.000 773.210 39.000 ;
        RECT 772.960 14.270 773.100 35.000 ;
        RECT 180.880 13.950 181.140 14.270 ;
        RECT 772.900 13.950 773.160 14.270 ;
        RECT 180.940 2.400 181.080 13.950 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 198.790 22.340 199.110 22.400 ;
        RECT 823.470 22.340 823.790 22.400 ;
        RECT 198.790 22.200 823.790 22.340 ;
        RECT 198.790 22.140 199.110 22.200 ;
        RECT 823.470 22.140 823.790 22.200 ;
      LAYER via ;
        RECT 198.820 22.140 199.080 22.400 ;
        RECT 823.500 22.140 823.760 22.400 ;
      LAYER met2 ;
        RECT 823.530 35.000 823.810 39.000 ;
        RECT 823.560 22.430 823.700 35.000 ;
        RECT 198.820 22.110 199.080 22.430 ;
        RECT 823.500 22.110 823.760 22.430 ;
        RECT 198.880 2.400 199.020 22.110 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 216.730 14.520 217.050 14.580 ;
        RECT 874.530 14.520 874.850 14.580 ;
        RECT 216.730 14.380 874.850 14.520 ;
        RECT 216.730 14.320 217.050 14.380 ;
        RECT 874.530 14.320 874.850 14.380 ;
      LAYER via ;
        RECT 216.760 14.320 217.020 14.580 ;
        RECT 874.560 14.320 874.820 14.580 ;
      LAYER met2 ;
        RECT 874.590 35.000 874.870 39.000 ;
        RECT 874.620 14.610 874.760 35.000 ;
        RECT 216.760 14.290 217.020 14.610 ;
        RECT 874.560 14.290 874.820 14.610 ;
        RECT 216.820 2.400 216.960 14.290 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 234.670 22.680 234.990 22.740 ;
        RECT 925.130 22.680 925.450 22.740 ;
        RECT 234.670 22.540 925.450 22.680 ;
        RECT 234.670 22.480 234.990 22.540 ;
        RECT 925.130 22.480 925.450 22.540 ;
      LAYER via ;
        RECT 234.700 22.480 234.960 22.740 ;
        RECT 925.160 22.480 925.420 22.740 ;
      LAYER met2 ;
        RECT 925.190 35.000 925.470 39.000 ;
        RECT 925.220 22.770 925.360 35.000 ;
        RECT 234.700 22.450 234.960 22.770 ;
        RECT 925.160 22.450 925.420 22.770 ;
        RECT 234.760 2.400 234.900 22.450 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.750 17.920 27.070 17.980 ;
        RECT 56.190 17.920 56.510 17.980 ;
        RECT 26.750 17.780 56.510 17.920 ;
        RECT 26.750 17.720 27.070 17.780 ;
        RECT 56.190 17.720 56.510 17.780 ;
      LAYER via ;
        RECT 26.780 17.720 27.040 17.980 ;
        RECT 56.220 17.720 56.480 17.980 ;
      LAYER met2 ;
        RECT 26.770 3277.755 27.050 3278.125 ;
        RECT 26.840 18.010 26.980 3277.755 ;
        RECT 26.780 17.690 27.040 18.010 ;
        RECT 56.220 17.690 56.480 18.010 ;
        RECT 56.280 2.400 56.420 17.690 ;
        RECT 56.070 -4.800 56.630 2.400 ;
      LAYER via2 ;
        RECT 26.770 3277.800 27.050 3278.080 ;
      LAYER met3 ;
        RECT 35.000 3279.320 39.000 3279.920 ;
        RECT 26.745 3278.090 27.075 3278.105 ;
        RECT 35.270 3278.090 35.570 3279.320 ;
        RECT 26.745 3277.790 35.570 3278.090 ;
        RECT 26.745 3277.775 27.075 3277.790 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 27.210 17.580 27.530 17.640 ;
        RECT 80.110 17.580 80.430 17.640 ;
        RECT 27.210 17.440 80.430 17.580 ;
        RECT 27.210 17.380 27.530 17.440 ;
        RECT 80.110 17.380 80.430 17.440 ;
      LAYER via ;
        RECT 27.240 17.380 27.500 17.640 ;
        RECT 80.140 17.380 80.400 17.640 ;
      LAYER met2 ;
        RECT 27.230 3381.795 27.510 3382.165 ;
        RECT 27.300 17.670 27.440 3381.795 ;
        RECT 27.240 17.350 27.500 17.670 ;
        RECT 80.140 17.350 80.400 17.670 ;
        RECT 80.200 2.400 80.340 17.350 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 27.230 3381.840 27.510 3382.120 ;
      LAYER met3 ;
        RECT 35.000 3382.680 39.000 3383.280 ;
        RECT 27.205 3382.130 27.535 3382.145 ;
        RECT 35.270 3382.130 35.570 3382.680 ;
        RECT 27.205 3381.830 35.570 3382.130 ;
        RECT 27.205 3381.815 27.535 3381.830 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.590 17.155 103.870 17.525 ;
        RECT 103.660 2.400 103.800 17.155 ;
        RECT 103.450 -4.800 104.010 2.400 ;
      LAYER via2 ;
        RECT 103.590 17.200 103.870 17.480 ;
      LAYER met3 ;
        RECT 2881.000 3252.120 2885.000 3252.720 ;
        RECT 2884.510 3250.210 2884.810 3252.120 ;
        RECT 2891.830 3250.210 2892.210 3250.220 ;
        RECT 2884.510 3249.910 2892.210 3250.210 ;
        RECT 2891.830 3249.900 2892.210 3249.910 ;
        RECT 103.565 17.490 103.895 17.505 ;
        RECT 2891.830 17.490 2892.210 17.500 ;
        RECT 103.565 17.190 2892.210 17.490 ;
        RECT 103.565 17.175 103.895 17.190 ;
        RECT 2891.830 17.180 2892.210 17.190 ;
      LAYER via3 ;
        RECT 2891.860 3249.900 2892.180 3250.220 ;
        RECT 2891.860 17.180 2892.180 17.500 ;
      LAYER met4 ;
        RECT 2891.855 3249.895 2892.185 3250.225 ;
        RECT 2891.870 17.505 2892.170 3249.895 ;
        RECT 2891.855 17.175 2892.185 17.505 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2831.850 3442.995 2832.130 3443.365 ;
        RECT 2831.920 3435.000 2832.060 3442.995 ;
        RECT 2831.890 3431.000 2832.170 3435.000 ;
        RECT 127.510 17.835 127.790 18.205 ;
        RECT 127.580 2.400 127.720 17.835 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 2831.850 3443.040 2832.130 3443.320 ;
        RECT 127.510 17.880 127.790 18.160 ;
      LAYER met3 ;
        RECT 2831.825 3443.330 2832.155 3443.345 ;
        RECT 2856.870 3443.330 2857.250 3443.340 ;
        RECT 2831.825 3443.030 2857.250 3443.330 ;
        RECT 2831.825 3443.015 2832.155 3443.030 ;
        RECT 2856.870 3443.020 2857.250 3443.030 ;
        RECT 127.485 18.170 127.815 18.185 ;
        RECT 2856.870 18.170 2857.250 18.180 ;
        RECT 127.485 17.870 2857.250 18.170 ;
        RECT 127.485 17.855 127.815 17.870 ;
        RECT 2856.870 17.860 2857.250 17.870 ;
      LAYER via3 ;
        RECT 2856.900 3443.020 2857.220 3443.340 ;
        RECT 2856.900 17.860 2857.220 18.180 ;
      LAYER met4 ;
        RECT 2856.895 3443.015 2857.225 3443.345 ;
        RECT 2856.910 18.185 2857.210 3443.015 ;
        RECT 2856.895 17.855 2857.225 18.185 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 16.475 26.590 16.845 ;
        RECT 26.380 2.400 26.520 16.475 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 26.310 16.520 26.590 16.800 ;
      LAYER met3 ;
        RECT 2890.910 3374.650 2891.290 3374.660 ;
        RECT 2884.510 3374.440 2891.290 3374.650 ;
        RECT 2881.000 3374.350 2891.290 3374.440 ;
        RECT 2881.000 3373.840 2885.000 3374.350 ;
        RECT 2890.910 3374.340 2891.290 3374.350 ;
        RECT 26.285 16.810 26.615 16.825 ;
        RECT 2890.910 16.810 2891.290 16.820 ;
        RECT 26.285 16.510 2891.290 16.810 ;
        RECT 26.285 16.495 26.615 16.510 ;
        RECT 2890.910 16.500 2891.290 16.510 ;
      LAYER via3 ;
        RECT 2890.940 3374.340 2891.260 3374.660 ;
        RECT 2890.940 16.500 2891.260 16.820 ;
      LAYER met4 ;
        RECT 2890.935 3374.335 2891.265 3374.665 ;
        RECT 2890.950 16.825 2891.250 3374.335 ;
        RECT 2890.935 16.495 2891.265 16.825 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2859.490 35.000 2859.770 39.000 ;
        RECT 2859.520 24.325 2859.660 35.000 ;
        RECT 32.290 23.955 32.570 24.325 ;
        RECT 2859.450 23.955 2859.730 24.325 ;
        RECT 32.360 2.400 32.500 23.955 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 32.290 24.000 32.570 24.280 ;
        RECT 2859.450 24.000 2859.730 24.280 ;
      LAYER met3 ;
        RECT 32.265 24.290 32.595 24.305 ;
        RECT 2859.425 24.290 2859.755 24.305 ;
        RECT 32.265 23.990 2859.755 24.290 ;
        RECT 32.265 23.975 32.595 23.990 ;
        RECT 2859.425 23.975 2859.755 23.990 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 117.120 -9.320 120.120 3529.000 ;
        RECT 877.120 -9.320 880.120 3529.000 ;
        RECT 1637.120 -9.320 1640.120 3529.000 ;
        RECT 2397.120 -9.320 2400.120 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 118.030 3523.010 119.210 3524.190 ;
        RECT 118.030 3521.410 119.210 3522.590 ;
        RECT 118.030 -2.910 119.210 -1.730 ;
        RECT 118.030 -4.510 119.210 -3.330 ;
        RECT 878.030 3523.010 879.210 3524.190 ;
        RECT 878.030 3521.410 879.210 3522.590 ;
        RECT 878.030 -2.910 879.210 -1.730 ;
        RECT 878.030 -4.510 879.210 -3.330 ;
        RECT 1638.030 3523.010 1639.210 3524.190 ;
        RECT 1638.030 3521.410 1639.210 3522.590 ;
        RECT 1638.030 -2.910 1639.210 -1.730 ;
        RECT 1638.030 -4.510 1639.210 -3.330 ;
        RECT 2398.030 3523.010 2399.210 3524.190 ;
        RECT 2398.030 3521.410 2399.210 3522.590 ;
        RECT 2398.030 -2.910 2399.210 -1.730 ;
        RECT 2398.030 -4.510 2399.210 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 117.120 3524.300 120.120 3524.310 ;
        RECT 877.120 3524.300 880.120 3524.310 ;
        RECT 1637.120 3524.300 1640.120 3524.310 ;
        RECT 2397.120 3524.300 2400.120 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 117.120 3521.290 120.120 3521.300 ;
        RECT 877.120 3521.290 880.120 3521.300 ;
        RECT 1637.120 3521.290 1640.120 3521.300 ;
        RECT 2397.120 3521.290 2400.120 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 117.120 -1.620 120.120 -1.610 ;
        RECT 877.120 -1.620 880.120 -1.610 ;
        RECT 1637.120 -1.620 1640.120 -1.610 ;
        RECT 2397.120 -1.620 2400.120 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 117.120 -4.630 120.120 -4.620 ;
        RECT 877.120 -4.630 880.120 -4.620 ;
        RECT 1637.120 -4.630 1640.120 -4.620 ;
        RECT 2397.120 -4.630 2400.120 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 497.120 -9.320 500.120 3529.000 ;
        RECT 1257.120 -9.320 1260.120 3529.000 ;
        RECT 2017.120 -9.320 2020.120 3529.000 ;
        RECT 2777.120 -9.320 2780.120 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 498.030 3527.710 499.210 3528.890 ;
        RECT 498.030 3526.110 499.210 3527.290 ;
        RECT 498.030 -7.610 499.210 -6.430 ;
        RECT 498.030 -9.210 499.210 -8.030 ;
        RECT 1258.030 3527.710 1259.210 3528.890 ;
        RECT 1258.030 3526.110 1259.210 3527.290 ;
        RECT 1258.030 -7.610 1259.210 -6.430 ;
        RECT 1258.030 -9.210 1259.210 -8.030 ;
        RECT 2018.030 3527.710 2019.210 3528.890 ;
        RECT 2018.030 3526.110 2019.210 3527.290 ;
        RECT 2018.030 -7.610 2019.210 -6.430 ;
        RECT 2018.030 -9.210 2019.210 -8.030 ;
        RECT 2778.030 3527.710 2779.210 3528.890 ;
        RECT 2778.030 3526.110 2779.210 3527.290 ;
        RECT 2778.030 -7.610 2779.210 -6.430 ;
        RECT 2778.030 -9.210 2779.210 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 497.120 3529.000 500.120 3529.010 ;
        RECT 1257.120 3529.000 1260.120 3529.010 ;
        RECT 2017.120 3529.000 2020.120 3529.010 ;
        RECT 2777.120 3529.000 2780.120 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 497.120 3525.990 500.120 3526.000 ;
        RECT 1257.120 3525.990 1260.120 3526.000 ;
        RECT 2017.120 3525.990 2020.120 3526.000 ;
        RECT 2777.120 3525.990 2780.120 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 497.120 -6.320 500.120 -6.310 ;
        RECT 1257.120 -6.320 1260.120 -6.310 ;
        RECT 2017.120 -6.320 2020.120 -6.310 ;
        RECT 2777.120 -6.320 2780.120 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 497.120 -9.330 500.120 -9.320 ;
        RECT 1257.120 -9.330 1260.120 -9.320 ;
        RECT 2017.120 -9.330 2020.120 -9.320 ;
        RECT 2777.120 -9.330 2780.120 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 40.520 45.795 2879.180 3424.205 ;
      LAYER met1 ;
        RECT 40.520 45.640 2879.180 3424.360 ;
      LAYER met2 ;
        RECT 48.780 3430.720 87.250 3431.000 ;
        RECT 88.090 3430.720 192.590 3431.000 ;
        RECT 193.430 3430.720 297.930 3431.000 ;
        RECT 298.770 3430.720 403.730 3431.000 ;
        RECT 404.570 3430.720 509.070 3431.000 ;
        RECT 509.910 3430.720 614.870 3431.000 ;
        RECT 615.710 3430.720 720.210 3431.000 ;
        RECT 721.050 3430.720 826.010 3431.000 ;
        RECT 826.850 3430.720 931.350 3431.000 ;
        RECT 932.190 3430.720 1037.150 3431.000 ;
        RECT 1037.990 3430.720 1142.490 3431.000 ;
        RECT 1143.330 3430.720 1248.290 3431.000 ;
        RECT 1249.130 3430.720 1353.630 3431.000 ;
        RECT 1354.470 3430.720 1459.430 3431.000 ;
        RECT 1460.270 3430.720 1564.770 3431.000 ;
        RECT 1565.610 3430.720 1670.570 3431.000 ;
        RECT 1671.410 3430.720 1775.910 3431.000 ;
        RECT 1776.750 3430.720 1881.710 3431.000 ;
        RECT 1882.550 3430.720 1987.050 3431.000 ;
        RECT 1987.890 3430.720 2092.850 3431.000 ;
        RECT 2093.690 3430.720 2198.190 3431.000 ;
        RECT 2199.030 3430.720 2303.990 3431.000 ;
        RECT 2304.830 3430.720 2409.330 3431.000 ;
        RECT 2410.170 3430.720 2515.130 3431.000 ;
        RECT 2515.970 3430.720 2620.470 3431.000 ;
        RECT 2621.310 3430.720 2726.270 3431.000 ;
        RECT 2727.110 3430.720 2831.610 3431.000 ;
        RECT 2832.450 3430.720 2870.810 3431.000 ;
        RECT 48.780 39.280 2870.810 3430.720 ;
        RECT 48.780 39.000 60.110 39.280 ;
        RECT 60.950 39.000 110.710 39.280 ;
        RECT 111.550 39.000 161.770 39.280 ;
        RECT 162.610 39.000 212.370 39.280 ;
        RECT 213.210 39.000 263.430 39.280 ;
        RECT 264.270 39.000 314.490 39.280 ;
        RECT 315.330 39.000 365.090 39.280 ;
        RECT 365.930 39.000 416.150 39.280 ;
        RECT 416.990 39.000 467.210 39.280 ;
        RECT 468.050 39.000 517.810 39.280 ;
        RECT 518.650 39.000 568.870 39.280 ;
        RECT 569.710 39.000 619.930 39.280 ;
        RECT 620.770 39.000 670.530 39.280 ;
        RECT 671.370 39.000 721.590 39.280 ;
        RECT 722.430 39.000 772.650 39.280 ;
        RECT 773.490 39.000 823.250 39.280 ;
        RECT 824.090 39.000 874.310 39.280 ;
        RECT 875.150 39.000 924.910 39.280 ;
        RECT 925.750 39.000 975.970 39.280 ;
        RECT 976.810 39.000 1027.030 39.280 ;
        RECT 1027.870 39.000 1077.630 39.280 ;
        RECT 1078.470 39.000 1128.690 39.280 ;
        RECT 1129.530 39.000 1179.750 39.280 ;
        RECT 1180.590 39.000 1230.350 39.280 ;
        RECT 1231.190 39.000 1281.410 39.280 ;
        RECT 1282.250 39.000 1332.470 39.280 ;
        RECT 1333.310 39.000 1383.070 39.280 ;
        RECT 1383.910 39.000 1434.130 39.280 ;
        RECT 1434.970 39.000 1485.190 39.280 ;
        RECT 1486.030 39.000 1535.790 39.280 ;
        RECT 1536.630 39.000 1586.850 39.280 ;
        RECT 1587.690 39.000 1637.450 39.280 ;
        RECT 1638.290 39.000 1688.510 39.280 ;
        RECT 1689.350 39.000 1739.570 39.280 ;
        RECT 1740.410 39.000 1790.170 39.280 ;
        RECT 1791.010 39.000 1841.230 39.280 ;
        RECT 1842.070 39.000 1892.290 39.280 ;
        RECT 1893.130 39.000 1942.890 39.280 ;
        RECT 1943.730 39.000 1993.950 39.280 ;
        RECT 1994.790 39.000 2045.010 39.280 ;
        RECT 2045.850 39.000 2095.610 39.280 ;
        RECT 2096.450 39.000 2146.670 39.280 ;
        RECT 2147.510 39.000 2197.730 39.280 ;
        RECT 2198.570 39.000 2248.330 39.280 ;
        RECT 2249.170 39.000 2299.390 39.280 ;
        RECT 2300.230 39.000 2349.990 39.280 ;
        RECT 2350.830 39.000 2401.050 39.280 ;
        RECT 2401.890 39.000 2452.110 39.280 ;
        RECT 2452.950 39.000 2502.710 39.280 ;
        RECT 2503.550 39.000 2553.770 39.280 ;
        RECT 2554.610 39.000 2604.830 39.280 ;
        RECT 2605.670 39.000 2655.430 39.280 ;
        RECT 2656.270 39.000 2706.490 39.280 ;
        RECT 2707.330 39.000 2757.550 39.280 ;
        RECT 2758.390 39.000 2808.150 39.280 ;
        RECT 2808.990 39.000 2859.210 39.280 ;
        RECT 2860.050 39.000 2870.810 39.280 ;
      LAYER met3 ;
        RECT 39.000 3383.680 2881.000 3424.285 ;
        RECT 39.400 3382.280 2881.000 3383.680 ;
        RECT 39.000 3374.840 2881.000 3382.280 ;
        RECT 39.000 3373.440 2880.600 3374.840 ;
        RECT 39.000 3280.320 2881.000 3373.440 ;
        RECT 39.400 3278.920 2881.000 3280.320 ;
        RECT 39.000 3253.120 2881.000 3278.920 ;
        RECT 39.000 3251.720 2880.600 3253.120 ;
        RECT 39.000 3177.640 2881.000 3251.720 ;
        RECT 39.400 3176.240 2881.000 3177.640 ;
        RECT 39.000 3132.080 2881.000 3176.240 ;
        RECT 39.000 3130.680 2880.600 3132.080 ;
        RECT 39.000 3074.280 2881.000 3130.680 ;
        RECT 39.400 3072.880 2881.000 3074.280 ;
        RECT 39.000 3010.360 2881.000 3072.880 ;
        RECT 39.000 3008.960 2880.600 3010.360 ;
        RECT 39.000 2971.600 2881.000 3008.960 ;
        RECT 39.400 2970.200 2881.000 2971.600 ;
        RECT 39.000 2889.320 2881.000 2970.200 ;
        RECT 39.000 2887.920 2880.600 2889.320 ;
        RECT 39.000 2868.240 2881.000 2887.920 ;
        RECT 39.400 2866.840 2881.000 2868.240 ;
        RECT 39.000 2767.600 2881.000 2866.840 ;
        RECT 39.000 2766.200 2880.600 2767.600 ;
        RECT 39.000 2765.560 2881.000 2766.200 ;
        RECT 39.400 2764.160 2881.000 2765.560 ;
        RECT 39.000 2662.200 2881.000 2764.160 ;
        RECT 39.400 2660.800 2881.000 2662.200 ;
        RECT 39.000 2646.560 2881.000 2660.800 ;
        RECT 39.000 2645.160 2880.600 2646.560 ;
        RECT 39.000 2559.520 2881.000 2645.160 ;
        RECT 39.400 2558.120 2881.000 2559.520 ;
        RECT 39.000 2524.840 2881.000 2558.120 ;
        RECT 39.000 2523.440 2880.600 2524.840 ;
        RECT 39.000 2456.160 2881.000 2523.440 ;
        RECT 39.400 2454.760 2881.000 2456.160 ;
        RECT 39.000 2403.120 2881.000 2454.760 ;
        RECT 39.000 2401.720 2880.600 2403.120 ;
        RECT 39.000 2353.480 2881.000 2401.720 ;
        RECT 39.400 2352.080 2881.000 2353.480 ;
        RECT 39.000 2282.080 2881.000 2352.080 ;
        RECT 39.000 2280.680 2880.600 2282.080 ;
        RECT 39.000 2250.120 2881.000 2280.680 ;
        RECT 39.400 2248.720 2881.000 2250.120 ;
        RECT 39.000 2160.360 2881.000 2248.720 ;
        RECT 39.000 2158.960 2880.600 2160.360 ;
        RECT 39.000 2147.440 2881.000 2158.960 ;
        RECT 39.400 2146.040 2881.000 2147.440 ;
        RECT 39.000 2044.080 2881.000 2146.040 ;
        RECT 39.400 2042.680 2881.000 2044.080 ;
        RECT 39.000 2039.320 2881.000 2042.680 ;
        RECT 39.000 2037.920 2880.600 2039.320 ;
        RECT 39.000 1941.400 2881.000 2037.920 ;
        RECT 39.400 1940.000 2881.000 1941.400 ;
        RECT 39.000 1917.600 2881.000 1940.000 ;
        RECT 39.000 1916.200 2880.600 1917.600 ;
        RECT 39.000 1838.040 2881.000 1916.200 ;
        RECT 39.400 1836.640 2881.000 1838.040 ;
        RECT 39.000 1796.560 2881.000 1836.640 ;
        RECT 39.000 1795.160 2880.600 1796.560 ;
        RECT 39.000 1735.360 2881.000 1795.160 ;
        RECT 39.400 1733.960 2881.000 1735.360 ;
        RECT 39.000 1674.840 2881.000 1733.960 ;
        RECT 39.000 1673.440 2880.600 1674.840 ;
        RECT 39.000 1632.000 2881.000 1673.440 ;
        RECT 39.400 1630.600 2881.000 1632.000 ;
        RECT 39.000 1553.120 2881.000 1630.600 ;
        RECT 39.000 1551.720 2880.600 1553.120 ;
        RECT 39.000 1529.320 2881.000 1551.720 ;
        RECT 39.400 1527.920 2881.000 1529.320 ;
        RECT 39.000 1432.080 2881.000 1527.920 ;
        RECT 39.000 1430.680 2880.600 1432.080 ;
        RECT 39.000 1425.960 2881.000 1430.680 ;
        RECT 39.400 1424.560 2881.000 1425.960 ;
        RECT 39.000 1323.280 2881.000 1424.560 ;
        RECT 39.400 1321.880 2881.000 1323.280 ;
        RECT 39.000 1310.360 2881.000 1321.880 ;
        RECT 39.000 1308.960 2880.600 1310.360 ;
        RECT 39.000 1219.920 2881.000 1308.960 ;
        RECT 39.400 1218.520 2881.000 1219.920 ;
        RECT 39.000 1189.320 2881.000 1218.520 ;
        RECT 39.000 1187.920 2880.600 1189.320 ;
        RECT 39.000 1117.240 2881.000 1187.920 ;
        RECT 39.400 1115.840 2881.000 1117.240 ;
        RECT 39.000 1067.600 2881.000 1115.840 ;
        RECT 39.000 1066.200 2880.600 1067.600 ;
        RECT 39.000 1013.880 2881.000 1066.200 ;
        RECT 39.400 1012.480 2881.000 1013.880 ;
        RECT 39.000 946.560 2881.000 1012.480 ;
        RECT 39.000 945.160 2880.600 946.560 ;
        RECT 39.000 911.200 2881.000 945.160 ;
        RECT 39.400 909.800 2881.000 911.200 ;
        RECT 39.000 824.840 2881.000 909.800 ;
        RECT 39.000 823.440 2880.600 824.840 ;
        RECT 39.000 807.840 2881.000 823.440 ;
        RECT 39.400 806.440 2881.000 807.840 ;
        RECT 39.000 705.160 2881.000 806.440 ;
        RECT 39.400 703.760 2881.000 705.160 ;
        RECT 39.000 703.120 2881.000 703.760 ;
        RECT 39.000 701.720 2880.600 703.120 ;
        RECT 39.000 601.800 2881.000 701.720 ;
        RECT 39.400 600.400 2881.000 601.800 ;
        RECT 39.000 582.080 2881.000 600.400 ;
        RECT 39.000 580.680 2880.600 582.080 ;
        RECT 39.000 499.120 2881.000 580.680 ;
        RECT 39.400 497.720 2881.000 499.120 ;
        RECT 39.000 460.360 2881.000 497.720 ;
        RECT 39.000 458.960 2880.600 460.360 ;
        RECT 39.000 395.760 2881.000 458.960 ;
        RECT 39.400 394.360 2881.000 395.760 ;
        RECT 39.000 339.320 2881.000 394.360 ;
        RECT 39.000 337.920 2880.600 339.320 ;
        RECT 39.000 293.080 2881.000 337.920 ;
        RECT 39.400 291.680 2881.000 293.080 ;
        RECT 39.000 217.600 2881.000 291.680 ;
        RECT 39.000 216.200 2880.600 217.600 ;
        RECT 39.000 189.720 2881.000 216.200 ;
        RECT 39.400 188.320 2881.000 189.720 ;
        RECT 39.000 96.560 2881.000 188.320 ;
        RECT 39.000 95.160 2880.600 96.560 ;
        RECT 39.000 87.040 2881.000 95.160 ;
        RECT 39.400 85.640 2881.000 87.040 ;
        RECT 39.000 45.715 2881.000 85.640 ;
      LAYER met4 ;
        RECT 48.720 45.640 117.120 3424.360 ;
        RECT 120.120 45.640 497.120 3424.360 ;
        RECT 500.120 45.640 877.120 3424.360 ;
        RECT 880.120 45.640 1257.120 3424.360 ;
        RECT 1260.120 45.640 1637.120 3424.360 ;
        RECT 1640.120 45.640 2017.120 3424.360 ;
        RECT 2020.120 45.640 2397.120 3424.360 ;
        RECT 2400.120 45.640 2777.120 3424.360 ;
        RECT 2780.120 45.640 2848.505 3424.360 ;
      LAYER met5 ;
        RECT 40.520 138.080 2879.180 3394.755 ;
      LAYER met5 ;
        RECT 40.520 99.785 2879.180 101.385 ;
        RECT 40.520 61.490 2879.180 63.090 ;
  END
END user_project_wrapper
END LIBRARY

